module SbufferData(
  input         clock,
  input         reset,
  input         io_writeReq_0_valid,
  input  [15:0] io_writeReq_0_bits_wvec,
  input  [7:0]  io_writeReq_0_bits_mask,
  input  [63:0] io_writeReq_0_bits_data,
  input  [32:0] io_writeReq_0_bits_wordOffset,
  input         io_writeReq_0_bits_wline,
  input         io_writeReq_1_valid,
  input  [15:0] io_writeReq_1_bits_wvec,
  input  [7:0]  io_writeReq_1_bits_mask,
  input  [63:0] io_writeReq_1_bits_data,
  input  [32:0] io_writeReq_1_bits_wordOffset,
  input         io_writeReq_1_bits_wline,
  input         io_maskFlushReq_0_valid,
  input  [15:0] io_maskFlushReq_0_bits_wvec,
  input         io_maskFlushReq_1_valid,
  input  [15:0] io_maskFlushReq_1_bits_wvec,
  output [7:0]  io_dataOut_0_0_0,
  output [7:0]  io_dataOut_0_0_1,
  output [7:0]  io_dataOut_0_0_2,
  output [7:0]  io_dataOut_0_0_3,
  output [7:0]  io_dataOut_0_0_4,
  output [7:0]  io_dataOut_0_0_5,
  output [7:0]  io_dataOut_0_0_6,
  output [7:0]  io_dataOut_0_0_7,
  output [7:0]  io_dataOut_0_1_0,
  output [7:0]  io_dataOut_0_1_1,
  output [7:0]  io_dataOut_0_1_2,
  output [7:0]  io_dataOut_0_1_3,
  output [7:0]  io_dataOut_0_1_4,
  output [7:0]  io_dataOut_0_1_5,
  output [7:0]  io_dataOut_0_1_6,
  output [7:0]  io_dataOut_0_1_7,
  output [7:0]  io_dataOut_0_2_0,
  output [7:0]  io_dataOut_0_2_1,
  output [7:0]  io_dataOut_0_2_2,
  output [7:0]  io_dataOut_0_2_3,
  output [7:0]  io_dataOut_0_2_4,
  output [7:0]  io_dataOut_0_2_5,
  output [7:0]  io_dataOut_0_2_6,
  output [7:0]  io_dataOut_0_2_7,
  output [7:0]  io_dataOut_0_3_0,
  output [7:0]  io_dataOut_0_3_1,
  output [7:0]  io_dataOut_0_3_2,
  output [7:0]  io_dataOut_0_3_3,
  output [7:0]  io_dataOut_0_3_4,
  output [7:0]  io_dataOut_0_3_5,
  output [7:0]  io_dataOut_0_3_6,
  output [7:0]  io_dataOut_0_3_7,
  output [7:0]  io_dataOut_0_4_0,
  output [7:0]  io_dataOut_0_4_1,
  output [7:0]  io_dataOut_0_4_2,
  output [7:0]  io_dataOut_0_4_3,
  output [7:0]  io_dataOut_0_4_4,
  output [7:0]  io_dataOut_0_4_5,
  output [7:0]  io_dataOut_0_4_6,
  output [7:0]  io_dataOut_0_4_7,
  output [7:0]  io_dataOut_0_5_0,
  output [7:0]  io_dataOut_0_5_1,
  output [7:0]  io_dataOut_0_5_2,
  output [7:0]  io_dataOut_0_5_3,
  output [7:0]  io_dataOut_0_5_4,
  output [7:0]  io_dataOut_0_5_5,
  output [7:0]  io_dataOut_0_5_6,
  output [7:0]  io_dataOut_0_5_7,
  output [7:0]  io_dataOut_0_6_0,
  output [7:0]  io_dataOut_0_6_1,
  output [7:0]  io_dataOut_0_6_2,
  output [7:0]  io_dataOut_0_6_3,
  output [7:0]  io_dataOut_0_6_4,
  output [7:0]  io_dataOut_0_6_5,
  output [7:0]  io_dataOut_0_6_6,
  output [7:0]  io_dataOut_0_6_7,
  output [7:0]  io_dataOut_0_7_0,
  output [7:0]  io_dataOut_0_7_1,
  output [7:0]  io_dataOut_0_7_2,
  output [7:0]  io_dataOut_0_7_3,
  output [7:0]  io_dataOut_0_7_4,
  output [7:0]  io_dataOut_0_7_5,
  output [7:0]  io_dataOut_0_7_6,
  output [7:0]  io_dataOut_0_7_7,
  output [7:0]  io_dataOut_1_0_0,
  output [7:0]  io_dataOut_1_0_1,
  output [7:0]  io_dataOut_1_0_2,
  output [7:0]  io_dataOut_1_0_3,
  output [7:0]  io_dataOut_1_0_4,
  output [7:0]  io_dataOut_1_0_5,
  output [7:0]  io_dataOut_1_0_6,
  output [7:0]  io_dataOut_1_0_7,
  output [7:0]  io_dataOut_1_1_0,
  output [7:0]  io_dataOut_1_1_1,
  output [7:0]  io_dataOut_1_1_2,
  output [7:0]  io_dataOut_1_1_3,
  output [7:0]  io_dataOut_1_1_4,
  output [7:0]  io_dataOut_1_1_5,
  output [7:0]  io_dataOut_1_1_6,
  output [7:0]  io_dataOut_1_1_7,
  output [7:0]  io_dataOut_1_2_0,
  output [7:0]  io_dataOut_1_2_1,
  output [7:0]  io_dataOut_1_2_2,
  output [7:0]  io_dataOut_1_2_3,
  output [7:0]  io_dataOut_1_2_4,
  output [7:0]  io_dataOut_1_2_5,
  output [7:0]  io_dataOut_1_2_6,
  output [7:0]  io_dataOut_1_2_7,
  output [7:0]  io_dataOut_1_3_0,
  output [7:0]  io_dataOut_1_3_1,
  output [7:0]  io_dataOut_1_3_2,
  output [7:0]  io_dataOut_1_3_3,
  output [7:0]  io_dataOut_1_3_4,
  output [7:0]  io_dataOut_1_3_5,
  output [7:0]  io_dataOut_1_3_6,
  output [7:0]  io_dataOut_1_3_7,
  output [7:0]  io_dataOut_1_4_0,
  output [7:0]  io_dataOut_1_4_1,
  output [7:0]  io_dataOut_1_4_2,
  output [7:0]  io_dataOut_1_4_3,
  output [7:0]  io_dataOut_1_4_4,
  output [7:0]  io_dataOut_1_4_5,
  output [7:0]  io_dataOut_1_4_6,
  output [7:0]  io_dataOut_1_4_7,
  output [7:0]  io_dataOut_1_5_0,
  output [7:0]  io_dataOut_1_5_1,
  output [7:0]  io_dataOut_1_5_2,
  output [7:0]  io_dataOut_1_5_3,
  output [7:0]  io_dataOut_1_5_4,
  output [7:0]  io_dataOut_1_5_5,
  output [7:0]  io_dataOut_1_5_6,
  output [7:0]  io_dataOut_1_5_7,
  output [7:0]  io_dataOut_1_6_0,
  output [7:0]  io_dataOut_1_6_1,
  output [7:0]  io_dataOut_1_6_2,
  output [7:0]  io_dataOut_1_6_3,
  output [7:0]  io_dataOut_1_6_4,
  output [7:0]  io_dataOut_1_6_5,
  output [7:0]  io_dataOut_1_6_6,
  output [7:0]  io_dataOut_1_6_7,
  output [7:0]  io_dataOut_1_7_0,
  output [7:0]  io_dataOut_1_7_1,
  output [7:0]  io_dataOut_1_7_2,
  output [7:0]  io_dataOut_1_7_3,
  output [7:0]  io_dataOut_1_7_4,
  output [7:0]  io_dataOut_1_7_5,
  output [7:0]  io_dataOut_1_7_6,
  output [7:0]  io_dataOut_1_7_7,
  output [7:0]  io_dataOut_2_0_0,
  output [7:0]  io_dataOut_2_0_1,
  output [7:0]  io_dataOut_2_0_2,
  output [7:0]  io_dataOut_2_0_3,
  output [7:0]  io_dataOut_2_0_4,
  output [7:0]  io_dataOut_2_0_5,
  output [7:0]  io_dataOut_2_0_6,
  output [7:0]  io_dataOut_2_0_7,
  output [7:0]  io_dataOut_2_1_0,
  output [7:0]  io_dataOut_2_1_1,
  output [7:0]  io_dataOut_2_1_2,
  output [7:0]  io_dataOut_2_1_3,
  output [7:0]  io_dataOut_2_1_4,
  output [7:0]  io_dataOut_2_1_5,
  output [7:0]  io_dataOut_2_1_6,
  output [7:0]  io_dataOut_2_1_7,
  output [7:0]  io_dataOut_2_2_0,
  output [7:0]  io_dataOut_2_2_1,
  output [7:0]  io_dataOut_2_2_2,
  output [7:0]  io_dataOut_2_2_3,
  output [7:0]  io_dataOut_2_2_4,
  output [7:0]  io_dataOut_2_2_5,
  output [7:0]  io_dataOut_2_2_6,
  output [7:0]  io_dataOut_2_2_7,
  output [7:0]  io_dataOut_2_3_0,
  output [7:0]  io_dataOut_2_3_1,
  output [7:0]  io_dataOut_2_3_2,
  output [7:0]  io_dataOut_2_3_3,
  output [7:0]  io_dataOut_2_3_4,
  output [7:0]  io_dataOut_2_3_5,
  output [7:0]  io_dataOut_2_3_6,
  output [7:0]  io_dataOut_2_3_7,
  output [7:0]  io_dataOut_2_4_0,
  output [7:0]  io_dataOut_2_4_1,
  output [7:0]  io_dataOut_2_4_2,
  output [7:0]  io_dataOut_2_4_3,
  output [7:0]  io_dataOut_2_4_4,
  output [7:0]  io_dataOut_2_4_5,
  output [7:0]  io_dataOut_2_4_6,
  output [7:0]  io_dataOut_2_4_7,
  output [7:0]  io_dataOut_2_5_0,
  output [7:0]  io_dataOut_2_5_1,
  output [7:0]  io_dataOut_2_5_2,
  output [7:0]  io_dataOut_2_5_3,
  output [7:0]  io_dataOut_2_5_4,
  output [7:0]  io_dataOut_2_5_5,
  output [7:0]  io_dataOut_2_5_6,
  output [7:0]  io_dataOut_2_5_7,
  output [7:0]  io_dataOut_2_6_0,
  output [7:0]  io_dataOut_2_6_1,
  output [7:0]  io_dataOut_2_6_2,
  output [7:0]  io_dataOut_2_6_3,
  output [7:0]  io_dataOut_2_6_4,
  output [7:0]  io_dataOut_2_6_5,
  output [7:0]  io_dataOut_2_6_6,
  output [7:0]  io_dataOut_2_6_7,
  output [7:0]  io_dataOut_2_7_0,
  output [7:0]  io_dataOut_2_7_1,
  output [7:0]  io_dataOut_2_7_2,
  output [7:0]  io_dataOut_2_7_3,
  output [7:0]  io_dataOut_2_7_4,
  output [7:0]  io_dataOut_2_7_5,
  output [7:0]  io_dataOut_2_7_6,
  output [7:0]  io_dataOut_2_7_7,
  output [7:0]  io_dataOut_3_0_0,
  output [7:0]  io_dataOut_3_0_1,
  output [7:0]  io_dataOut_3_0_2,
  output [7:0]  io_dataOut_3_0_3,
  output [7:0]  io_dataOut_3_0_4,
  output [7:0]  io_dataOut_3_0_5,
  output [7:0]  io_dataOut_3_0_6,
  output [7:0]  io_dataOut_3_0_7,
  output [7:0]  io_dataOut_3_1_0,
  output [7:0]  io_dataOut_3_1_1,
  output [7:0]  io_dataOut_3_1_2,
  output [7:0]  io_dataOut_3_1_3,
  output [7:0]  io_dataOut_3_1_4,
  output [7:0]  io_dataOut_3_1_5,
  output [7:0]  io_dataOut_3_1_6,
  output [7:0]  io_dataOut_3_1_7,
  output [7:0]  io_dataOut_3_2_0,
  output [7:0]  io_dataOut_3_2_1,
  output [7:0]  io_dataOut_3_2_2,
  output [7:0]  io_dataOut_3_2_3,
  output [7:0]  io_dataOut_3_2_4,
  output [7:0]  io_dataOut_3_2_5,
  output [7:0]  io_dataOut_3_2_6,
  output [7:0]  io_dataOut_3_2_7,
  output [7:0]  io_dataOut_3_3_0,
  output [7:0]  io_dataOut_3_3_1,
  output [7:0]  io_dataOut_3_3_2,
  output [7:0]  io_dataOut_3_3_3,
  output [7:0]  io_dataOut_3_3_4,
  output [7:0]  io_dataOut_3_3_5,
  output [7:0]  io_dataOut_3_3_6,
  output [7:0]  io_dataOut_3_3_7,
  output [7:0]  io_dataOut_3_4_0,
  output [7:0]  io_dataOut_3_4_1,
  output [7:0]  io_dataOut_3_4_2,
  output [7:0]  io_dataOut_3_4_3,
  output [7:0]  io_dataOut_3_4_4,
  output [7:0]  io_dataOut_3_4_5,
  output [7:0]  io_dataOut_3_4_6,
  output [7:0]  io_dataOut_3_4_7,
  output [7:0]  io_dataOut_3_5_0,
  output [7:0]  io_dataOut_3_5_1,
  output [7:0]  io_dataOut_3_5_2,
  output [7:0]  io_dataOut_3_5_3,
  output [7:0]  io_dataOut_3_5_4,
  output [7:0]  io_dataOut_3_5_5,
  output [7:0]  io_dataOut_3_5_6,
  output [7:0]  io_dataOut_3_5_7,
  output [7:0]  io_dataOut_3_6_0,
  output [7:0]  io_dataOut_3_6_1,
  output [7:0]  io_dataOut_3_6_2,
  output [7:0]  io_dataOut_3_6_3,
  output [7:0]  io_dataOut_3_6_4,
  output [7:0]  io_dataOut_3_6_5,
  output [7:0]  io_dataOut_3_6_6,
  output [7:0]  io_dataOut_3_6_7,
  output [7:0]  io_dataOut_3_7_0,
  output [7:0]  io_dataOut_3_7_1,
  output [7:0]  io_dataOut_3_7_2,
  output [7:0]  io_dataOut_3_7_3,
  output [7:0]  io_dataOut_3_7_4,
  output [7:0]  io_dataOut_3_7_5,
  output [7:0]  io_dataOut_3_7_6,
  output [7:0]  io_dataOut_3_7_7,
  output [7:0]  io_dataOut_4_0_0,
  output [7:0]  io_dataOut_4_0_1,
  output [7:0]  io_dataOut_4_0_2,
  output [7:0]  io_dataOut_4_0_3,
  output [7:0]  io_dataOut_4_0_4,
  output [7:0]  io_dataOut_4_0_5,
  output [7:0]  io_dataOut_4_0_6,
  output [7:0]  io_dataOut_4_0_7,
  output [7:0]  io_dataOut_4_1_0,
  output [7:0]  io_dataOut_4_1_1,
  output [7:0]  io_dataOut_4_1_2,
  output [7:0]  io_dataOut_4_1_3,
  output [7:0]  io_dataOut_4_1_4,
  output [7:0]  io_dataOut_4_1_5,
  output [7:0]  io_dataOut_4_1_6,
  output [7:0]  io_dataOut_4_1_7,
  output [7:0]  io_dataOut_4_2_0,
  output [7:0]  io_dataOut_4_2_1,
  output [7:0]  io_dataOut_4_2_2,
  output [7:0]  io_dataOut_4_2_3,
  output [7:0]  io_dataOut_4_2_4,
  output [7:0]  io_dataOut_4_2_5,
  output [7:0]  io_dataOut_4_2_6,
  output [7:0]  io_dataOut_4_2_7,
  output [7:0]  io_dataOut_4_3_0,
  output [7:0]  io_dataOut_4_3_1,
  output [7:0]  io_dataOut_4_3_2,
  output [7:0]  io_dataOut_4_3_3,
  output [7:0]  io_dataOut_4_3_4,
  output [7:0]  io_dataOut_4_3_5,
  output [7:0]  io_dataOut_4_3_6,
  output [7:0]  io_dataOut_4_3_7,
  output [7:0]  io_dataOut_4_4_0,
  output [7:0]  io_dataOut_4_4_1,
  output [7:0]  io_dataOut_4_4_2,
  output [7:0]  io_dataOut_4_4_3,
  output [7:0]  io_dataOut_4_4_4,
  output [7:0]  io_dataOut_4_4_5,
  output [7:0]  io_dataOut_4_4_6,
  output [7:0]  io_dataOut_4_4_7,
  output [7:0]  io_dataOut_4_5_0,
  output [7:0]  io_dataOut_4_5_1,
  output [7:0]  io_dataOut_4_5_2,
  output [7:0]  io_dataOut_4_5_3,
  output [7:0]  io_dataOut_4_5_4,
  output [7:0]  io_dataOut_4_5_5,
  output [7:0]  io_dataOut_4_5_6,
  output [7:0]  io_dataOut_4_5_7,
  output [7:0]  io_dataOut_4_6_0,
  output [7:0]  io_dataOut_4_6_1,
  output [7:0]  io_dataOut_4_6_2,
  output [7:0]  io_dataOut_4_6_3,
  output [7:0]  io_dataOut_4_6_4,
  output [7:0]  io_dataOut_4_6_5,
  output [7:0]  io_dataOut_4_6_6,
  output [7:0]  io_dataOut_4_6_7,
  output [7:0]  io_dataOut_4_7_0,
  output [7:0]  io_dataOut_4_7_1,
  output [7:0]  io_dataOut_4_7_2,
  output [7:0]  io_dataOut_4_7_3,
  output [7:0]  io_dataOut_4_7_4,
  output [7:0]  io_dataOut_4_7_5,
  output [7:0]  io_dataOut_4_7_6,
  output [7:0]  io_dataOut_4_7_7,
  output [7:0]  io_dataOut_5_0_0,
  output [7:0]  io_dataOut_5_0_1,
  output [7:0]  io_dataOut_5_0_2,
  output [7:0]  io_dataOut_5_0_3,
  output [7:0]  io_dataOut_5_0_4,
  output [7:0]  io_dataOut_5_0_5,
  output [7:0]  io_dataOut_5_0_6,
  output [7:0]  io_dataOut_5_0_7,
  output [7:0]  io_dataOut_5_1_0,
  output [7:0]  io_dataOut_5_1_1,
  output [7:0]  io_dataOut_5_1_2,
  output [7:0]  io_dataOut_5_1_3,
  output [7:0]  io_dataOut_5_1_4,
  output [7:0]  io_dataOut_5_1_5,
  output [7:0]  io_dataOut_5_1_6,
  output [7:0]  io_dataOut_5_1_7,
  output [7:0]  io_dataOut_5_2_0,
  output [7:0]  io_dataOut_5_2_1,
  output [7:0]  io_dataOut_5_2_2,
  output [7:0]  io_dataOut_5_2_3,
  output [7:0]  io_dataOut_5_2_4,
  output [7:0]  io_dataOut_5_2_5,
  output [7:0]  io_dataOut_5_2_6,
  output [7:0]  io_dataOut_5_2_7,
  output [7:0]  io_dataOut_5_3_0,
  output [7:0]  io_dataOut_5_3_1,
  output [7:0]  io_dataOut_5_3_2,
  output [7:0]  io_dataOut_5_3_3,
  output [7:0]  io_dataOut_5_3_4,
  output [7:0]  io_dataOut_5_3_5,
  output [7:0]  io_dataOut_5_3_6,
  output [7:0]  io_dataOut_5_3_7,
  output [7:0]  io_dataOut_5_4_0,
  output [7:0]  io_dataOut_5_4_1,
  output [7:0]  io_dataOut_5_4_2,
  output [7:0]  io_dataOut_5_4_3,
  output [7:0]  io_dataOut_5_4_4,
  output [7:0]  io_dataOut_5_4_5,
  output [7:0]  io_dataOut_5_4_6,
  output [7:0]  io_dataOut_5_4_7,
  output [7:0]  io_dataOut_5_5_0,
  output [7:0]  io_dataOut_5_5_1,
  output [7:0]  io_dataOut_5_5_2,
  output [7:0]  io_dataOut_5_5_3,
  output [7:0]  io_dataOut_5_5_4,
  output [7:0]  io_dataOut_5_5_5,
  output [7:0]  io_dataOut_5_5_6,
  output [7:0]  io_dataOut_5_5_7,
  output [7:0]  io_dataOut_5_6_0,
  output [7:0]  io_dataOut_5_6_1,
  output [7:0]  io_dataOut_5_6_2,
  output [7:0]  io_dataOut_5_6_3,
  output [7:0]  io_dataOut_5_6_4,
  output [7:0]  io_dataOut_5_6_5,
  output [7:0]  io_dataOut_5_6_6,
  output [7:0]  io_dataOut_5_6_7,
  output [7:0]  io_dataOut_5_7_0,
  output [7:0]  io_dataOut_5_7_1,
  output [7:0]  io_dataOut_5_7_2,
  output [7:0]  io_dataOut_5_7_3,
  output [7:0]  io_dataOut_5_7_4,
  output [7:0]  io_dataOut_5_7_5,
  output [7:0]  io_dataOut_5_7_6,
  output [7:0]  io_dataOut_5_7_7,
  output [7:0]  io_dataOut_6_0_0,
  output [7:0]  io_dataOut_6_0_1,
  output [7:0]  io_dataOut_6_0_2,
  output [7:0]  io_dataOut_6_0_3,
  output [7:0]  io_dataOut_6_0_4,
  output [7:0]  io_dataOut_6_0_5,
  output [7:0]  io_dataOut_6_0_6,
  output [7:0]  io_dataOut_6_0_7,
  output [7:0]  io_dataOut_6_1_0,
  output [7:0]  io_dataOut_6_1_1,
  output [7:0]  io_dataOut_6_1_2,
  output [7:0]  io_dataOut_6_1_3,
  output [7:0]  io_dataOut_6_1_4,
  output [7:0]  io_dataOut_6_1_5,
  output [7:0]  io_dataOut_6_1_6,
  output [7:0]  io_dataOut_6_1_7,
  output [7:0]  io_dataOut_6_2_0,
  output [7:0]  io_dataOut_6_2_1,
  output [7:0]  io_dataOut_6_2_2,
  output [7:0]  io_dataOut_6_2_3,
  output [7:0]  io_dataOut_6_2_4,
  output [7:0]  io_dataOut_6_2_5,
  output [7:0]  io_dataOut_6_2_6,
  output [7:0]  io_dataOut_6_2_7,
  output [7:0]  io_dataOut_6_3_0,
  output [7:0]  io_dataOut_6_3_1,
  output [7:0]  io_dataOut_6_3_2,
  output [7:0]  io_dataOut_6_3_3,
  output [7:0]  io_dataOut_6_3_4,
  output [7:0]  io_dataOut_6_3_5,
  output [7:0]  io_dataOut_6_3_6,
  output [7:0]  io_dataOut_6_3_7,
  output [7:0]  io_dataOut_6_4_0,
  output [7:0]  io_dataOut_6_4_1,
  output [7:0]  io_dataOut_6_4_2,
  output [7:0]  io_dataOut_6_4_3,
  output [7:0]  io_dataOut_6_4_4,
  output [7:0]  io_dataOut_6_4_5,
  output [7:0]  io_dataOut_6_4_6,
  output [7:0]  io_dataOut_6_4_7,
  output [7:0]  io_dataOut_6_5_0,
  output [7:0]  io_dataOut_6_5_1,
  output [7:0]  io_dataOut_6_5_2,
  output [7:0]  io_dataOut_6_5_3,
  output [7:0]  io_dataOut_6_5_4,
  output [7:0]  io_dataOut_6_5_5,
  output [7:0]  io_dataOut_6_5_6,
  output [7:0]  io_dataOut_6_5_7,
  output [7:0]  io_dataOut_6_6_0,
  output [7:0]  io_dataOut_6_6_1,
  output [7:0]  io_dataOut_6_6_2,
  output [7:0]  io_dataOut_6_6_3,
  output [7:0]  io_dataOut_6_6_4,
  output [7:0]  io_dataOut_6_6_5,
  output [7:0]  io_dataOut_6_6_6,
  output [7:0]  io_dataOut_6_6_7,
  output [7:0]  io_dataOut_6_7_0,
  output [7:0]  io_dataOut_6_7_1,
  output [7:0]  io_dataOut_6_7_2,
  output [7:0]  io_dataOut_6_7_3,
  output [7:0]  io_dataOut_6_7_4,
  output [7:0]  io_dataOut_6_7_5,
  output [7:0]  io_dataOut_6_7_6,
  output [7:0]  io_dataOut_6_7_7,
  output [7:0]  io_dataOut_7_0_0,
  output [7:0]  io_dataOut_7_0_1,
  output [7:0]  io_dataOut_7_0_2,
  output [7:0]  io_dataOut_7_0_3,
  output [7:0]  io_dataOut_7_0_4,
  output [7:0]  io_dataOut_7_0_5,
  output [7:0]  io_dataOut_7_0_6,
  output [7:0]  io_dataOut_7_0_7,
  output [7:0]  io_dataOut_7_1_0,
  output [7:0]  io_dataOut_7_1_1,
  output [7:0]  io_dataOut_7_1_2,
  output [7:0]  io_dataOut_7_1_3,
  output [7:0]  io_dataOut_7_1_4,
  output [7:0]  io_dataOut_7_1_5,
  output [7:0]  io_dataOut_7_1_6,
  output [7:0]  io_dataOut_7_1_7,
  output [7:0]  io_dataOut_7_2_0,
  output [7:0]  io_dataOut_7_2_1,
  output [7:0]  io_dataOut_7_2_2,
  output [7:0]  io_dataOut_7_2_3,
  output [7:0]  io_dataOut_7_2_4,
  output [7:0]  io_dataOut_7_2_5,
  output [7:0]  io_dataOut_7_2_6,
  output [7:0]  io_dataOut_7_2_7,
  output [7:0]  io_dataOut_7_3_0,
  output [7:0]  io_dataOut_7_3_1,
  output [7:0]  io_dataOut_7_3_2,
  output [7:0]  io_dataOut_7_3_3,
  output [7:0]  io_dataOut_7_3_4,
  output [7:0]  io_dataOut_7_3_5,
  output [7:0]  io_dataOut_7_3_6,
  output [7:0]  io_dataOut_7_3_7,
  output [7:0]  io_dataOut_7_4_0,
  output [7:0]  io_dataOut_7_4_1,
  output [7:0]  io_dataOut_7_4_2,
  output [7:0]  io_dataOut_7_4_3,
  output [7:0]  io_dataOut_7_4_4,
  output [7:0]  io_dataOut_7_4_5,
  output [7:0]  io_dataOut_7_4_6,
  output [7:0]  io_dataOut_7_4_7,
  output [7:0]  io_dataOut_7_5_0,
  output [7:0]  io_dataOut_7_5_1,
  output [7:0]  io_dataOut_7_5_2,
  output [7:0]  io_dataOut_7_5_3,
  output [7:0]  io_dataOut_7_5_4,
  output [7:0]  io_dataOut_7_5_5,
  output [7:0]  io_dataOut_7_5_6,
  output [7:0]  io_dataOut_7_5_7,
  output [7:0]  io_dataOut_7_6_0,
  output [7:0]  io_dataOut_7_6_1,
  output [7:0]  io_dataOut_7_6_2,
  output [7:0]  io_dataOut_7_6_3,
  output [7:0]  io_dataOut_7_6_4,
  output [7:0]  io_dataOut_7_6_5,
  output [7:0]  io_dataOut_7_6_6,
  output [7:0]  io_dataOut_7_6_7,
  output [7:0]  io_dataOut_7_7_0,
  output [7:0]  io_dataOut_7_7_1,
  output [7:0]  io_dataOut_7_7_2,
  output [7:0]  io_dataOut_7_7_3,
  output [7:0]  io_dataOut_7_7_4,
  output [7:0]  io_dataOut_7_7_5,
  output [7:0]  io_dataOut_7_7_6,
  output [7:0]  io_dataOut_7_7_7,
  output [7:0]  io_dataOut_8_0_0,
  output [7:0]  io_dataOut_8_0_1,
  output [7:0]  io_dataOut_8_0_2,
  output [7:0]  io_dataOut_8_0_3,
  output [7:0]  io_dataOut_8_0_4,
  output [7:0]  io_dataOut_8_0_5,
  output [7:0]  io_dataOut_8_0_6,
  output [7:0]  io_dataOut_8_0_7,
  output [7:0]  io_dataOut_8_1_0,
  output [7:0]  io_dataOut_8_1_1,
  output [7:0]  io_dataOut_8_1_2,
  output [7:0]  io_dataOut_8_1_3,
  output [7:0]  io_dataOut_8_1_4,
  output [7:0]  io_dataOut_8_1_5,
  output [7:0]  io_dataOut_8_1_6,
  output [7:0]  io_dataOut_8_1_7,
  output [7:0]  io_dataOut_8_2_0,
  output [7:0]  io_dataOut_8_2_1,
  output [7:0]  io_dataOut_8_2_2,
  output [7:0]  io_dataOut_8_2_3,
  output [7:0]  io_dataOut_8_2_4,
  output [7:0]  io_dataOut_8_2_5,
  output [7:0]  io_dataOut_8_2_6,
  output [7:0]  io_dataOut_8_2_7,
  output [7:0]  io_dataOut_8_3_0,
  output [7:0]  io_dataOut_8_3_1,
  output [7:0]  io_dataOut_8_3_2,
  output [7:0]  io_dataOut_8_3_3,
  output [7:0]  io_dataOut_8_3_4,
  output [7:0]  io_dataOut_8_3_5,
  output [7:0]  io_dataOut_8_3_6,
  output [7:0]  io_dataOut_8_3_7,
  output [7:0]  io_dataOut_8_4_0,
  output [7:0]  io_dataOut_8_4_1,
  output [7:0]  io_dataOut_8_4_2,
  output [7:0]  io_dataOut_8_4_3,
  output [7:0]  io_dataOut_8_4_4,
  output [7:0]  io_dataOut_8_4_5,
  output [7:0]  io_dataOut_8_4_6,
  output [7:0]  io_dataOut_8_4_7,
  output [7:0]  io_dataOut_8_5_0,
  output [7:0]  io_dataOut_8_5_1,
  output [7:0]  io_dataOut_8_5_2,
  output [7:0]  io_dataOut_8_5_3,
  output [7:0]  io_dataOut_8_5_4,
  output [7:0]  io_dataOut_8_5_5,
  output [7:0]  io_dataOut_8_5_6,
  output [7:0]  io_dataOut_8_5_7,
  output [7:0]  io_dataOut_8_6_0,
  output [7:0]  io_dataOut_8_6_1,
  output [7:0]  io_dataOut_8_6_2,
  output [7:0]  io_dataOut_8_6_3,
  output [7:0]  io_dataOut_8_6_4,
  output [7:0]  io_dataOut_8_6_5,
  output [7:0]  io_dataOut_8_6_6,
  output [7:0]  io_dataOut_8_6_7,
  output [7:0]  io_dataOut_8_7_0,
  output [7:0]  io_dataOut_8_7_1,
  output [7:0]  io_dataOut_8_7_2,
  output [7:0]  io_dataOut_8_7_3,
  output [7:0]  io_dataOut_8_7_4,
  output [7:0]  io_dataOut_8_7_5,
  output [7:0]  io_dataOut_8_7_6,
  output [7:0]  io_dataOut_8_7_7,
  output [7:0]  io_dataOut_9_0_0,
  output [7:0]  io_dataOut_9_0_1,
  output [7:0]  io_dataOut_9_0_2,
  output [7:0]  io_dataOut_9_0_3,
  output [7:0]  io_dataOut_9_0_4,
  output [7:0]  io_dataOut_9_0_5,
  output [7:0]  io_dataOut_9_0_6,
  output [7:0]  io_dataOut_9_0_7,
  output [7:0]  io_dataOut_9_1_0,
  output [7:0]  io_dataOut_9_1_1,
  output [7:0]  io_dataOut_9_1_2,
  output [7:0]  io_dataOut_9_1_3,
  output [7:0]  io_dataOut_9_1_4,
  output [7:0]  io_dataOut_9_1_5,
  output [7:0]  io_dataOut_9_1_6,
  output [7:0]  io_dataOut_9_1_7,
  output [7:0]  io_dataOut_9_2_0,
  output [7:0]  io_dataOut_9_2_1,
  output [7:0]  io_dataOut_9_2_2,
  output [7:0]  io_dataOut_9_2_3,
  output [7:0]  io_dataOut_9_2_4,
  output [7:0]  io_dataOut_9_2_5,
  output [7:0]  io_dataOut_9_2_6,
  output [7:0]  io_dataOut_9_2_7,
  output [7:0]  io_dataOut_9_3_0,
  output [7:0]  io_dataOut_9_3_1,
  output [7:0]  io_dataOut_9_3_2,
  output [7:0]  io_dataOut_9_3_3,
  output [7:0]  io_dataOut_9_3_4,
  output [7:0]  io_dataOut_9_3_5,
  output [7:0]  io_dataOut_9_3_6,
  output [7:0]  io_dataOut_9_3_7,
  output [7:0]  io_dataOut_9_4_0,
  output [7:0]  io_dataOut_9_4_1,
  output [7:0]  io_dataOut_9_4_2,
  output [7:0]  io_dataOut_9_4_3,
  output [7:0]  io_dataOut_9_4_4,
  output [7:0]  io_dataOut_9_4_5,
  output [7:0]  io_dataOut_9_4_6,
  output [7:0]  io_dataOut_9_4_7,
  output [7:0]  io_dataOut_9_5_0,
  output [7:0]  io_dataOut_9_5_1,
  output [7:0]  io_dataOut_9_5_2,
  output [7:0]  io_dataOut_9_5_3,
  output [7:0]  io_dataOut_9_5_4,
  output [7:0]  io_dataOut_9_5_5,
  output [7:0]  io_dataOut_9_5_6,
  output [7:0]  io_dataOut_9_5_7,
  output [7:0]  io_dataOut_9_6_0,
  output [7:0]  io_dataOut_9_6_1,
  output [7:0]  io_dataOut_9_6_2,
  output [7:0]  io_dataOut_9_6_3,
  output [7:0]  io_dataOut_9_6_4,
  output [7:0]  io_dataOut_9_6_5,
  output [7:0]  io_dataOut_9_6_6,
  output [7:0]  io_dataOut_9_6_7,
  output [7:0]  io_dataOut_9_7_0,
  output [7:0]  io_dataOut_9_7_1,
  output [7:0]  io_dataOut_9_7_2,
  output [7:0]  io_dataOut_9_7_3,
  output [7:0]  io_dataOut_9_7_4,
  output [7:0]  io_dataOut_9_7_5,
  output [7:0]  io_dataOut_9_7_6,
  output [7:0]  io_dataOut_9_7_7,
  output [7:0]  io_dataOut_10_0_0,
  output [7:0]  io_dataOut_10_0_1,
  output [7:0]  io_dataOut_10_0_2,
  output [7:0]  io_dataOut_10_0_3,
  output [7:0]  io_dataOut_10_0_4,
  output [7:0]  io_dataOut_10_0_5,
  output [7:0]  io_dataOut_10_0_6,
  output [7:0]  io_dataOut_10_0_7,
  output [7:0]  io_dataOut_10_1_0,
  output [7:0]  io_dataOut_10_1_1,
  output [7:0]  io_dataOut_10_1_2,
  output [7:0]  io_dataOut_10_1_3,
  output [7:0]  io_dataOut_10_1_4,
  output [7:0]  io_dataOut_10_1_5,
  output [7:0]  io_dataOut_10_1_6,
  output [7:0]  io_dataOut_10_1_7,
  output [7:0]  io_dataOut_10_2_0,
  output [7:0]  io_dataOut_10_2_1,
  output [7:0]  io_dataOut_10_2_2,
  output [7:0]  io_dataOut_10_2_3,
  output [7:0]  io_dataOut_10_2_4,
  output [7:0]  io_dataOut_10_2_5,
  output [7:0]  io_dataOut_10_2_6,
  output [7:0]  io_dataOut_10_2_7,
  output [7:0]  io_dataOut_10_3_0,
  output [7:0]  io_dataOut_10_3_1,
  output [7:0]  io_dataOut_10_3_2,
  output [7:0]  io_dataOut_10_3_3,
  output [7:0]  io_dataOut_10_3_4,
  output [7:0]  io_dataOut_10_3_5,
  output [7:0]  io_dataOut_10_3_6,
  output [7:0]  io_dataOut_10_3_7,
  output [7:0]  io_dataOut_10_4_0,
  output [7:0]  io_dataOut_10_4_1,
  output [7:0]  io_dataOut_10_4_2,
  output [7:0]  io_dataOut_10_4_3,
  output [7:0]  io_dataOut_10_4_4,
  output [7:0]  io_dataOut_10_4_5,
  output [7:0]  io_dataOut_10_4_6,
  output [7:0]  io_dataOut_10_4_7,
  output [7:0]  io_dataOut_10_5_0,
  output [7:0]  io_dataOut_10_5_1,
  output [7:0]  io_dataOut_10_5_2,
  output [7:0]  io_dataOut_10_5_3,
  output [7:0]  io_dataOut_10_5_4,
  output [7:0]  io_dataOut_10_5_5,
  output [7:0]  io_dataOut_10_5_6,
  output [7:0]  io_dataOut_10_5_7,
  output [7:0]  io_dataOut_10_6_0,
  output [7:0]  io_dataOut_10_6_1,
  output [7:0]  io_dataOut_10_6_2,
  output [7:0]  io_dataOut_10_6_3,
  output [7:0]  io_dataOut_10_6_4,
  output [7:0]  io_dataOut_10_6_5,
  output [7:0]  io_dataOut_10_6_6,
  output [7:0]  io_dataOut_10_6_7,
  output [7:0]  io_dataOut_10_7_0,
  output [7:0]  io_dataOut_10_7_1,
  output [7:0]  io_dataOut_10_7_2,
  output [7:0]  io_dataOut_10_7_3,
  output [7:0]  io_dataOut_10_7_4,
  output [7:0]  io_dataOut_10_7_5,
  output [7:0]  io_dataOut_10_7_6,
  output [7:0]  io_dataOut_10_7_7,
  output [7:0]  io_dataOut_11_0_0,
  output [7:0]  io_dataOut_11_0_1,
  output [7:0]  io_dataOut_11_0_2,
  output [7:0]  io_dataOut_11_0_3,
  output [7:0]  io_dataOut_11_0_4,
  output [7:0]  io_dataOut_11_0_5,
  output [7:0]  io_dataOut_11_0_6,
  output [7:0]  io_dataOut_11_0_7,
  output [7:0]  io_dataOut_11_1_0,
  output [7:0]  io_dataOut_11_1_1,
  output [7:0]  io_dataOut_11_1_2,
  output [7:0]  io_dataOut_11_1_3,
  output [7:0]  io_dataOut_11_1_4,
  output [7:0]  io_dataOut_11_1_5,
  output [7:0]  io_dataOut_11_1_6,
  output [7:0]  io_dataOut_11_1_7,
  output [7:0]  io_dataOut_11_2_0,
  output [7:0]  io_dataOut_11_2_1,
  output [7:0]  io_dataOut_11_2_2,
  output [7:0]  io_dataOut_11_2_3,
  output [7:0]  io_dataOut_11_2_4,
  output [7:0]  io_dataOut_11_2_5,
  output [7:0]  io_dataOut_11_2_6,
  output [7:0]  io_dataOut_11_2_7,
  output [7:0]  io_dataOut_11_3_0,
  output [7:0]  io_dataOut_11_3_1,
  output [7:0]  io_dataOut_11_3_2,
  output [7:0]  io_dataOut_11_3_3,
  output [7:0]  io_dataOut_11_3_4,
  output [7:0]  io_dataOut_11_3_5,
  output [7:0]  io_dataOut_11_3_6,
  output [7:0]  io_dataOut_11_3_7,
  output [7:0]  io_dataOut_11_4_0,
  output [7:0]  io_dataOut_11_4_1,
  output [7:0]  io_dataOut_11_4_2,
  output [7:0]  io_dataOut_11_4_3,
  output [7:0]  io_dataOut_11_4_4,
  output [7:0]  io_dataOut_11_4_5,
  output [7:0]  io_dataOut_11_4_6,
  output [7:0]  io_dataOut_11_4_7,
  output [7:0]  io_dataOut_11_5_0,
  output [7:0]  io_dataOut_11_5_1,
  output [7:0]  io_dataOut_11_5_2,
  output [7:0]  io_dataOut_11_5_3,
  output [7:0]  io_dataOut_11_5_4,
  output [7:0]  io_dataOut_11_5_5,
  output [7:0]  io_dataOut_11_5_6,
  output [7:0]  io_dataOut_11_5_7,
  output [7:0]  io_dataOut_11_6_0,
  output [7:0]  io_dataOut_11_6_1,
  output [7:0]  io_dataOut_11_6_2,
  output [7:0]  io_dataOut_11_6_3,
  output [7:0]  io_dataOut_11_6_4,
  output [7:0]  io_dataOut_11_6_5,
  output [7:0]  io_dataOut_11_6_6,
  output [7:0]  io_dataOut_11_6_7,
  output [7:0]  io_dataOut_11_7_0,
  output [7:0]  io_dataOut_11_7_1,
  output [7:0]  io_dataOut_11_7_2,
  output [7:0]  io_dataOut_11_7_3,
  output [7:0]  io_dataOut_11_7_4,
  output [7:0]  io_dataOut_11_7_5,
  output [7:0]  io_dataOut_11_7_6,
  output [7:0]  io_dataOut_11_7_7,
  output [7:0]  io_dataOut_12_0_0,
  output [7:0]  io_dataOut_12_0_1,
  output [7:0]  io_dataOut_12_0_2,
  output [7:0]  io_dataOut_12_0_3,
  output [7:0]  io_dataOut_12_0_4,
  output [7:0]  io_dataOut_12_0_5,
  output [7:0]  io_dataOut_12_0_6,
  output [7:0]  io_dataOut_12_0_7,
  output [7:0]  io_dataOut_12_1_0,
  output [7:0]  io_dataOut_12_1_1,
  output [7:0]  io_dataOut_12_1_2,
  output [7:0]  io_dataOut_12_1_3,
  output [7:0]  io_dataOut_12_1_4,
  output [7:0]  io_dataOut_12_1_5,
  output [7:0]  io_dataOut_12_1_6,
  output [7:0]  io_dataOut_12_1_7,
  output [7:0]  io_dataOut_12_2_0,
  output [7:0]  io_dataOut_12_2_1,
  output [7:0]  io_dataOut_12_2_2,
  output [7:0]  io_dataOut_12_2_3,
  output [7:0]  io_dataOut_12_2_4,
  output [7:0]  io_dataOut_12_2_5,
  output [7:0]  io_dataOut_12_2_6,
  output [7:0]  io_dataOut_12_2_7,
  output [7:0]  io_dataOut_12_3_0,
  output [7:0]  io_dataOut_12_3_1,
  output [7:0]  io_dataOut_12_3_2,
  output [7:0]  io_dataOut_12_3_3,
  output [7:0]  io_dataOut_12_3_4,
  output [7:0]  io_dataOut_12_3_5,
  output [7:0]  io_dataOut_12_3_6,
  output [7:0]  io_dataOut_12_3_7,
  output [7:0]  io_dataOut_12_4_0,
  output [7:0]  io_dataOut_12_4_1,
  output [7:0]  io_dataOut_12_4_2,
  output [7:0]  io_dataOut_12_4_3,
  output [7:0]  io_dataOut_12_4_4,
  output [7:0]  io_dataOut_12_4_5,
  output [7:0]  io_dataOut_12_4_6,
  output [7:0]  io_dataOut_12_4_7,
  output [7:0]  io_dataOut_12_5_0,
  output [7:0]  io_dataOut_12_5_1,
  output [7:0]  io_dataOut_12_5_2,
  output [7:0]  io_dataOut_12_5_3,
  output [7:0]  io_dataOut_12_5_4,
  output [7:0]  io_dataOut_12_5_5,
  output [7:0]  io_dataOut_12_5_6,
  output [7:0]  io_dataOut_12_5_7,
  output [7:0]  io_dataOut_12_6_0,
  output [7:0]  io_dataOut_12_6_1,
  output [7:0]  io_dataOut_12_6_2,
  output [7:0]  io_dataOut_12_6_3,
  output [7:0]  io_dataOut_12_6_4,
  output [7:0]  io_dataOut_12_6_5,
  output [7:0]  io_dataOut_12_6_6,
  output [7:0]  io_dataOut_12_6_7,
  output [7:0]  io_dataOut_12_7_0,
  output [7:0]  io_dataOut_12_7_1,
  output [7:0]  io_dataOut_12_7_2,
  output [7:0]  io_dataOut_12_7_3,
  output [7:0]  io_dataOut_12_7_4,
  output [7:0]  io_dataOut_12_7_5,
  output [7:0]  io_dataOut_12_7_6,
  output [7:0]  io_dataOut_12_7_7,
  output [7:0]  io_dataOut_13_0_0,
  output [7:0]  io_dataOut_13_0_1,
  output [7:0]  io_dataOut_13_0_2,
  output [7:0]  io_dataOut_13_0_3,
  output [7:0]  io_dataOut_13_0_4,
  output [7:0]  io_dataOut_13_0_5,
  output [7:0]  io_dataOut_13_0_6,
  output [7:0]  io_dataOut_13_0_7,
  output [7:0]  io_dataOut_13_1_0,
  output [7:0]  io_dataOut_13_1_1,
  output [7:0]  io_dataOut_13_1_2,
  output [7:0]  io_dataOut_13_1_3,
  output [7:0]  io_dataOut_13_1_4,
  output [7:0]  io_dataOut_13_1_5,
  output [7:0]  io_dataOut_13_1_6,
  output [7:0]  io_dataOut_13_1_7,
  output [7:0]  io_dataOut_13_2_0,
  output [7:0]  io_dataOut_13_2_1,
  output [7:0]  io_dataOut_13_2_2,
  output [7:0]  io_dataOut_13_2_3,
  output [7:0]  io_dataOut_13_2_4,
  output [7:0]  io_dataOut_13_2_5,
  output [7:0]  io_dataOut_13_2_6,
  output [7:0]  io_dataOut_13_2_7,
  output [7:0]  io_dataOut_13_3_0,
  output [7:0]  io_dataOut_13_3_1,
  output [7:0]  io_dataOut_13_3_2,
  output [7:0]  io_dataOut_13_3_3,
  output [7:0]  io_dataOut_13_3_4,
  output [7:0]  io_dataOut_13_3_5,
  output [7:0]  io_dataOut_13_3_6,
  output [7:0]  io_dataOut_13_3_7,
  output [7:0]  io_dataOut_13_4_0,
  output [7:0]  io_dataOut_13_4_1,
  output [7:0]  io_dataOut_13_4_2,
  output [7:0]  io_dataOut_13_4_3,
  output [7:0]  io_dataOut_13_4_4,
  output [7:0]  io_dataOut_13_4_5,
  output [7:0]  io_dataOut_13_4_6,
  output [7:0]  io_dataOut_13_4_7,
  output [7:0]  io_dataOut_13_5_0,
  output [7:0]  io_dataOut_13_5_1,
  output [7:0]  io_dataOut_13_5_2,
  output [7:0]  io_dataOut_13_5_3,
  output [7:0]  io_dataOut_13_5_4,
  output [7:0]  io_dataOut_13_5_5,
  output [7:0]  io_dataOut_13_5_6,
  output [7:0]  io_dataOut_13_5_7,
  output [7:0]  io_dataOut_13_6_0,
  output [7:0]  io_dataOut_13_6_1,
  output [7:0]  io_dataOut_13_6_2,
  output [7:0]  io_dataOut_13_6_3,
  output [7:0]  io_dataOut_13_6_4,
  output [7:0]  io_dataOut_13_6_5,
  output [7:0]  io_dataOut_13_6_6,
  output [7:0]  io_dataOut_13_6_7,
  output [7:0]  io_dataOut_13_7_0,
  output [7:0]  io_dataOut_13_7_1,
  output [7:0]  io_dataOut_13_7_2,
  output [7:0]  io_dataOut_13_7_3,
  output [7:0]  io_dataOut_13_7_4,
  output [7:0]  io_dataOut_13_7_5,
  output [7:0]  io_dataOut_13_7_6,
  output [7:0]  io_dataOut_13_7_7,
  output [7:0]  io_dataOut_14_0_0,
  output [7:0]  io_dataOut_14_0_1,
  output [7:0]  io_dataOut_14_0_2,
  output [7:0]  io_dataOut_14_0_3,
  output [7:0]  io_dataOut_14_0_4,
  output [7:0]  io_dataOut_14_0_5,
  output [7:0]  io_dataOut_14_0_6,
  output [7:0]  io_dataOut_14_0_7,
  output [7:0]  io_dataOut_14_1_0,
  output [7:0]  io_dataOut_14_1_1,
  output [7:0]  io_dataOut_14_1_2,
  output [7:0]  io_dataOut_14_1_3,
  output [7:0]  io_dataOut_14_1_4,
  output [7:0]  io_dataOut_14_1_5,
  output [7:0]  io_dataOut_14_1_6,
  output [7:0]  io_dataOut_14_1_7,
  output [7:0]  io_dataOut_14_2_0,
  output [7:0]  io_dataOut_14_2_1,
  output [7:0]  io_dataOut_14_2_2,
  output [7:0]  io_dataOut_14_2_3,
  output [7:0]  io_dataOut_14_2_4,
  output [7:0]  io_dataOut_14_2_5,
  output [7:0]  io_dataOut_14_2_6,
  output [7:0]  io_dataOut_14_2_7,
  output [7:0]  io_dataOut_14_3_0,
  output [7:0]  io_dataOut_14_3_1,
  output [7:0]  io_dataOut_14_3_2,
  output [7:0]  io_dataOut_14_3_3,
  output [7:0]  io_dataOut_14_3_4,
  output [7:0]  io_dataOut_14_3_5,
  output [7:0]  io_dataOut_14_3_6,
  output [7:0]  io_dataOut_14_3_7,
  output [7:0]  io_dataOut_14_4_0,
  output [7:0]  io_dataOut_14_4_1,
  output [7:0]  io_dataOut_14_4_2,
  output [7:0]  io_dataOut_14_4_3,
  output [7:0]  io_dataOut_14_4_4,
  output [7:0]  io_dataOut_14_4_5,
  output [7:0]  io_dataOut_14_4_6,
  output [7:0]  io_dataOut_14_4_7,
  output [7:0]  io_dataOut_14_5_0,
  output [7:0]  io_dataOut_14_5_1,
  output [7:0]  io_dataOut_14_5_2,
  output [7:0]  io_dataOut_14_5_3,
  output [7:0]  io_dataOut_14_5_4,
  output [7:0]  io_dataOut_14_5_5,
  output [7:0]  io_dataOut_14_5_6,
  output [7:0]  io_dataOut_14_5_7,
  output [7:0]  io_dataOut_14_6_0,
  output [7:0]  io_dataOut_14_6_1,
  output [7:0]  io_dataOut_14_6_2,
  output [7:0]  io_dataOut_14_6_3,
  output [7:0]  io_dataOut_14_6_4,
  output [7:0]  io_dataOut_14_6_5,
  output [7:0]  io_dataOut_14_6_6,
  output [7:0]  io_dataOut_14_6_7,
  output [7:0]  io_dataOut_14_7_0,
  output [7:0]  io_dataOut_14_7_1,
  output [7:0]  io_dataOut_14_7_2,
  output [7:0]  io_dataOut_14_7_3,
  output [7:0]  io_dataOut_14_7_4,
  output [7:0]  io_dataOut_14_7_5,
  output [7:0]  io_dataOut_14_7_6,
  output [7:0]  io_dataOut_14_7_7,
  output [7:0]  io_dataOut_15_0_0,
  output [7:0]  io_dataOut_15_0_1,
  output [7:0]  io_dataOut_15_0_2,
  output [7:0]  io_dataOut_15_0_3,
  output [7:0]  io_dataOut_15_0_4,
  output [7:0]  io_dataOut_15_0_5,
  output [7:0]  io_dataOut_15_0_6,
  output [7:0]  io_dataOut_15_0_7,
  output [7:0]  io_dataOut_15_1_0,
  output [7:0]  io_dataOut_15_1_1,
  output [7:0]  io_dataOut_15_1_2,
  output [7:0]  io_dataOut_15_1_3,
  output [7:0]  io_dataOut_15_1_4,
  output [7:0]  io_dataOut_15_1_5,
  output [7:0]  io_dataOut_15_1_6,
  output [7:0]  io_dataOut_15_1_7,
  output [7:0]  io_dataOut_15_2_0,
  output [7:0]  io_dataOut_15_2_1,
  output [7:0]  io_dataOut_15_2_2,
  output [7:0]  io_dataOut_15_2_3,
  output [7:0]  io_dataOut_15_2_4,
  output [7:0]  io_dataOut_15_2_5,
  output [7:0]  io_dataOut_15_2_6,
  output [7:0]  io_dataOut_15_2_7,
  output [7:0]  io_dataOut_15_3_0,
  output [7:0]  io_dataOut_15_3_1,
  output [7:0]  io_dataOut_15_3_2,
  output [7:0]  io_dataOut_15_3_3,
  output [7:0]  io_dataOut_15_3_4,
  output [7:0]  io_dataOut_15_3_5,
  output [7:0]  io_dataOut_15_3_6,
  output [7:0]  io_dataOut_15_3_7,
  output [7:0]  io_dataOut_15_4_0,
  output [7:0]  io_dataOut_15_4_1,
  output [7:0]  io_dataOut_15_4_2,
  output [7:0]  io_dataOut_15_4_3,
  output [7:0]  io_dataOut_15_4_4,
  output [7:0]  io_dataOut_15_4_5,
  output [7:0]  io_dataOut_15_4_6,
  output [7:0]  io_dataOut_15_4_7,
  output [7:0]  io_dataOut_15_5_0,
  output [7:0]  io_dataOut_15_5_1,
  output [7:0]  io_dataOut_15_5_2,
  output [7:0]  io_dataOut_15_5_3,
  output [7:0]  io_dataOut_15_5_4,
  output [7:0]  io_dataOut_15_5_5,
  output [7:0]  io_dataOut_15_5_6,
  output [7:0]  io_dataOut_15_5_7,
  output [7:0]  io_dataOut_15_6_0,
  output [7:0]  io_dataOut_15_6_1,
  output [7:0]  io_dataOut_15_6_2,
  output [7:0]  io_dataOut_15_6_3,
  output [7:0]  io_dataOut_15_6_4,
  output [7:0]  io_dataOut_15_6_5,
  output [7:0]  io_dataOut_15_6_6,
  output [7:0]  io_dataOut_15_6_7,
  output [7:0]  io_dataOut_15_7_0,
  output [7:0]  io_dataOut_15_7_1,
  output [7:0]  io_dataOut_15_7_2,
  output [7:0]  io_dataOut_15_7_3,
  output [7:0]  io_dataOut_15_7_4,
  output [7:0]  io_dataOut_15_7_5,
  output [7:0]  io_dataOut_15_7_6,
  output [7:0]  io_dataOut_15_7_7,
  output        io_maskOut_0_0_0,
  output        io_maskOut_0_0_1,
  output        io_maskOut_0_0_2,
  output        io_maskOut_0_0_3,
  output        io_maskOut_0_0_4,
  output        io_maskOut_0_0_5,
  output        io_maskOut_0_0_6,
  output        io_maskOut_0_0_7,
  output        io_maskOut_0_1_0,
  output        io_maskOut_0_1_1,
  output        io_maskOut_0_1_2,
  output        io_maskOut_0_1_3,
  output        io_maskOut_0_1_4,
  output        io_maskOut_0_1_5,
  output        io_maskOut_0_1_6,
  output        io_maskOut_0_1_7,
  output        io_maskOut_0_2_0,
  output        io_maskOut_0_2_1,
  output        io_maskOut_0_2_2,
  output        io_maskOut_0_2_3,
  output        io_maskOut_0_2_4,
  output        io_maskOut_0_2_5,
  output        io_maskOut_0_2_6,
  output        io_maskOut_0_2_7,
  output        io_maskOut_0_3_0,
  output        io_maskOut_0_3_1,
  output        io_maskOut_0_3_2,
  output        io_maskOut_0_3_3,
  output        io_maskOut_0_3_4,
  output        io_maskOut_0_3_5,
  output        io_maskOut_0_3_6,
  output        io_maskOut_0_3_7,
  output        io_maskOut_0_4_0,
  output        io_maskOut_0_4_1,
  output        io_maskOut_0_4_2,
  output        io_maskOut_0_4_3,
  output        io_maskOut_0_4_4,
  output        io_maskOut_0_4_5,
  output        io_maskOut_0_4_6,
  output        io_maskOut_0_4_7,
  output        io_maskOut_0_5_0,
  output        io_maskOut_0_5_1,
  output        io_maskOut_0_5_2,
  output        io_maskOut_0_5_3,
  output        io_maskOut_0_5_4,
  output        io_maskOut_0_5_5,
  output        io_maskOut_0_5_6,
  output        io_maskOut_0_5_7,
  output        io_maskOut_0_6_0,
  output        io_maskOut_0_6_1,
  output        io_maskOut_0_6_2,
  output        io_maskOut_0_6_3,
  output        io_maskOut_0_6_4,
  output        io_maskOut_0_6_5,
  output        io_maskOut_0_6_6,
  output        io_maskOut_0_6_7,
  output        io_maskOut_0_7_0,
  output        io_maskOut_0_7_1,
  output        io_maskOut_0_7_2,
  output        io_maskOut_0_7_3,
  output        io_maskOut_0_7_4,
  output        io_maskOut_0_7_5,
  output        io_maskOut_0_7_6,
  output        io_maskOut_0_7_7,
  output        io_maskOut_1_0_0,
  output        io_maskOut_1_0_1,
  output        io_maskOut_1_0_2,
  output        io_maskOut_1_0_3,
  output        io_maskOut_1_0_4,
  output        io_maskOut_1_0_5,
  output        io_maskOut_1_0_6,
  output        io_maskOut_1_0_7,
  output        io_maskOut_1_1_0,
  output        io_maskOut_1_1_1,
  output        io_maskOut_1_1_2,
  output        io_maskOut_1_1_3,
  output        io_maskOut_1_1_4,
  output        io_maskOut_1_1_5,
  output        io_maskOut_1_1_6,
  output        io_maskOut_1_1_7,
  output        io_maskOut_1_2_0,
  output        io_maskOut_1_2_1,
  output        io_maskOut_1_2_2,
  output        io_maskOut_1_2_3,
  output        io_maskOut_1_2_4,
  output        io_maskOut_1_2_5,
  output        io_maskOut_1_2_6,
  output        io_maskOut_1_2_7,
  output        io_maskOut_1_3_0,
  output        io_maskOut_1_3_1,
  output        io_maskOut_1_3_2,
  output        io_maskOut_1_3_3,
  output        io_maskOut_1_3_4,
  output        io_maskOut_1_3_5,
  output        io_maskOut_1_3_6,
  output        io_maskOut_1_3_7,
  output        io_maskOut_1_4_0,
  output        io_maskOut_1_4_1,
  output        io_maskOut_1_4_2,
  output        io_maskOut_1_4_3,
  output        io_maskOut_1_4_4,
  output        io_maskOut_1_4_5,
  output        io_maskOut_1_4_6,
  output        io_maskOut_1_4_7,
  output        io_maskOut_1_5_0,
  output        io_maskOut_1_5_1,
  output        io_maskOut_1_5_2,
  output        io_maskOut_1_5_3,
  output        io_maskOut_1_5_4,
  output        io_maskOut_1_5_5,
  output        io_maskOut_1_5_6,
  output        io_maskOut_1_5_7,
  output        io_maskOut_1_6_0,
  output        io_maskOut_1_6_1,
  output        io_maskOut_1_6_2,
  output        io_maskOut_1_6_3,
  output        io_maskOut_1_6_4,
  output        io_maskOut_1_6_5,
  output        io_maskOut_1_6_6,
  output        io_maskOut_1_6_7,
  output        io_maskOut_1_7_0,
  output        io_maskOut_1_7_1,
  output        io_maskOut_1_7_2,
  output        io_maskOut_1_7_3,
  output        io_maskOut_1_7_4,
  output        io_maskOut_1_7_5,
  output        io_maskOut_1_7_6,
  output        io_maskOut_1_7_7,
  output        io_maskOut_2_0_0,
  output        io_maskOut_2_0_1,
  output        io_maskOut_2_0_2,
  output        io_maskOut_2_0_3,
  output        io_maskOut_2_0_4,
  output        io_maskOut_2_0_5,
  output        io_maskOut_2_0_6,
  output        io_maskOut_2_0_7,
  output        io_maskOut_2_1_0,
  output        io_maskOut_2_1_1,
  output        io_maskOut_2_1_2,
  output        io_maskOut_2_1_3,
  output        io_maskOut_2_1_4,
  output        io_maskOut_2_1_5,
  output        io_maskOut_2_1_6,
  output        io_maskOut_2_1_7,
  output        io_maskOut_2_2_0,
  output        io_maskOut_2_2_1,
  output        io_maskOut_2_2_2,
  output        io_maskOut_2_2_3,
  output        io_maskOut_2_2_4,
  output        io_maskOut_2_2_5,
  output        io_maskOut_2_2_6,
  output        io_maskOut_2_2_7,
  output        io_maskOut_2_3_0,
  output        io_maskOut_2_3_1,
  output        io_maskOut_2_3_2,
  output        io_maskOut_2_3_3,
  output        io_maskOut_2_3_4,
  output        io_maskOut_2_3_5,
  output        io_maskOut_2_3_6,
  output        io_maskOut_2_3_7,
  output        io_maskOut_2_4_0,
  output        io_maskOut_2_4_1,
  output        io_maskOut_2_4_2,
  output        io_maskOut_2_4_3,
  output        io_maskOut_2_4_4,
  output        io_maskOut_2_4_5,
  output        io_maskOut_2_4_6,
  output        io_maskOut_2_4_7,
  output        io_maskOut_2_5_0,
  output        io_maskOut_2_5_1,
  output        io_maskOut_2_5_2,
  output        io_maskOut_2_5_3,
  output        io_maskOut_2_5_4,
  output        io_maskOut_2_5_5,
  output        io_maskOut_2_5_6,
  output        io_maskOut_2_5_7,
  output        io_maskOut_2_6_0,
  output        io_maskOut_2_6_1,
  output        io_maskOut_2_6_2,
  output        io_maskOut_2_6_3,
  output        io_maskOut_2_6_4,
  output        io_maskOut_2_6_5,
  output        io_maskOut_2_6_6,
  output        io_maskOut_2_6_7,
  output        io_maskOut_2_7_0,
  output        io_maskOut_2_7_1,
  output        io_maskOut_2_7_2,
  output        io_maskOut_2_7_3,
  output        io_maskOut_2_7_4,
  output        io_maskOut_2_7_5,
  output        io_maskOut_2_7_6,
  output        io_maskOut_2_7_7,
  output        io_maskOut_3_0_0,
  output        io_maskOut_3_0_1,
  output        io_maskOut_3_0_2,
  output        io_maskOut_3_0_3,
  output        io_maskOut_3_0_4,
  output        io_maskOut_3_0_5,
  output        io_maskOut_3_0_6,
  output        io_maskOut_3_0_7,
  output        io_maskOut_3_1_0,
  output        io_maskOut_3_1_1,
  output        io_maskOut_3_1_2,
  output        io_maskOut_3_1_3,
  output        io_maskOut_3_1_4,
  output        io_maskOut_3_1_5,
  output        io_maskOut_3_1_6,
  output        io_maskOut_3_1_7,
  output        io_maskOut_3_2_0,
  output        io_maskOut_3_2_1,
  output        io_maskOut_3_2_2,
  output        io_maskOut_3_2_3,
  output        io_maskOut_3_2_4,
  output        io_maskOut_3_2_5,
  output        io_maskOut_3_2_6,
  output        io_maskOut_3_2_7,
  output        io_maskOut_3_3_0,
  output        io_maskOut_3_3_1,
  output        io_maskOut_3_3_2,
  output        io_maskOut_3_3_3,
  output        io_maskOut_3_3_4,
  output        io_maskOut_3_3_5,
  output        io_maskOut_3_3_6,
  output        io_maskOut_3_3_7,
  output        io_maskOut_3_4_0,
  output        io_maskOut_3_4_1,
  output        io_maskOut_3_4_2,
  output        io_maskOut_3_4_3,
  output        io_maskOut_3_4_4,
  output        io_maskOut_3_4_5,
  output        io_maskOut_3_4_6,
  output        io_maskOut_3_4_7,
  output        io_maskOut_3_5_0,
  output        io_maskOut_3_5_1,
  output        io_maskOut_3_5_2,
  output        io_maskOut_3_5_3,
  output        io_maskOut_3_5_4,
  output        io_maskOut_3_5_5,
  output        io_maskOut_3_5_6,
  output        io_maskOut_3_5_7,
  output        io_maskOut_3_6_0,
  output        io_maskOut_3_6_1,
  output        io_maskOut_3_6_2,
  output        io_maskOut_3_6_3,
  output        io_maskOut_3_6_4,
  output        io_maskOut_3_6_5,
  output        io_maskOut_3_6_6,
  output        io_maskOut_3_6_7,
  output        io_maskOut_3_7_0,
  output        io_maskOut_3_7_1,
  output        io_maskOut_3_7_2,
  output        io_maskOut_3_7_3,
  output        io_maskOut_3_7_4,
  output        io_maskOut_3_7_5,
  output        io_maskOut_3_7_6,
  output        io_maskOut_3_7_7,
  output        io_maskOut_4_0_0,
  output        io_maskOut_4_0_1,
  output        io_maskOut_4_0_2,
  output        io_maskOut_4_0_3,
  output        io_maskOut_4_0_4,
  output        io_maskOut_4_0_5,
  output        io_maskOut_4_0_6,
  output        io_maskOut_4_0_7,
  output        io_maskOut_4_1_0,
  output        io_maskOut_4_1_1,
  output        io_maskOut_4_1_2,
  output        io_maskOut_4_1_3,
  output        io_maskOut_4_1_4,
  output        io_maskOut_4_1_5,
  output        io_maskOut_4_1_6,
  output        io_maskOut_4_1_7,
  output        io_maskOut_4_2_0,
  output        io_maskOut_4_2_1,
  output        io_maskOut_4_2_2,
  output        io_maskOut_4_2_3,
  output        io_maskOut_4_2_4,
  output        io_maskOut_4_2_5,
  output        io_maskOut_4_2_6,
  output        io_maskOut_4_2_7,
  output        io_maskOut_4_3_0,
  output        io_maskOut_4_3_1,
  output        io_maskOut_4_3_2,
  output        io_maskOut_4_3_3,
  output        io_maskOut_4_3_4,
  output        io_maskOut_4_3_5,
  output        io_maskOut_4_3_6,
  output        io_maskOut_4_3_7,
  output        io_maskOut_4_4_0,
  output        io_maskOut_4_4_1,
  output        io_maskOut_4_4_2,
  output        io_maskOut_4_4_3,
  output        io_maskOut_4_4_4,
  output        io_maskOut_4_4_5,
  output        io_maskOut_4_4_6,
  output        io_maskOut_4_4_7,
  output        io_maskOut_4_5_0,
  output        io_maskOut_4_5_1,
  output        io_maskOut_4_5_2,
  output        io_maskOut_4_5_3,
  output        io_maskOut_4_5_4,
  output        io_maskOut_4_5_5,
  output        io_maskOut_4_5_6,
  output        io_maskOut_4_5_7,
  output        io_maskOut_4_6_0,
  output        io_maskOut_4_6_1,
  output        io_maskOut_4_6_2,
  output        io_maskOut_4_6_3,
  output        io_maskOut_4_6_4,
  output        io_maskOut_4_6_5,
  output        io_maskOut_4_6_6,
  output        io_maskOut_4_6_7,
  output        io_maskOut_4_7_0,
  output        io_maskOut_4_7_1,
  output        io_maskOut_4_7_2,
  output        io_maskOut_4_7_3,
  output        io_maskOut_4_7_4,
  output        io_maskOut_4_7_5,
  output        io_maskOut_4_7_6,
  output        io_maskOut_4_7_7,
  output        io_maskOut_5_0_0,
  output        io_maskOut_5_0_1,
  output        io_maskOut_5_0_2,
  output        io_maskOut_5_0_3,
  output        io_maskOut_5_0_4,
  output        io_maskOut_5_0_5,
  output        io_maskOut_5_0_6,
  output        io_maskOut_5_0_7,
  output        io_maskOut_5_1_0,
  output        io_maskOut_5_1_1,
  output        io_maskOut_5_1_2,
  output        io_maskOut_5_1_3,
  output        io_maskOut_5_1_4,
  output        io_maskOut_5_1_5,
  output        io_maskOut_5_1_6,
  output        io_maskOut_5_1_7,
  output        io_maskOut_5_2_0,
  output        io_maskOut_5_2_1,
  output        io_maskOut_5_2_2,
  output        io_maskOut_5_2_3,
  output        io_maskOut_5_2_4,
  output        io_maskOut_5_2_5,
  output        io_maskOut_5_2_6,
  output        io_maskOut_5_2_7,
  output        io_maskOut_5_3_0,
  output        io_maskOut_5_3_1,
  output        io_maskOut_5_3_2,
  output        io_maskOut_5_3_3,
  output        io_maskOut_5_3_4,
  output        io_maskOut_5_3_5,
  output        io_maskOut_5_3_6,
  output        io_maskOut_5_3_7,
  output        io_maskOut_5_4_0,
  output        io_maskOut_5_4_1,
  output        io_maskOut_5_4_2,
  output        io_maskOut_5_4_3,
  output        io_maskOut_5_4_4,
  output        io_maskOut_5_4_5,
  output        io_maskOut_5_4_6,
  output        io_maskOut_5_4_7,
  output        io_maskOut_5_5_0,
  output        io_maskOut_5_5_1,
  output        io_maskOut_5_5_2,
  output        io_maskOut_5_5_3,
  output        io_maskOut_5_5_4,
  output        io_maskOut_5_5_5,
  output        io_maskOut_5_5_6,
  output        io_maskOut_5_5_7,
  output        io_maskOut_5_6_0,
  output        io_maskOut_5_6_1,
  output        io_maskOut_5_6_2,
  output        io_maskOut_5_6_3,
  output        io_maskOut_5_6_4,
  output        io_maskOut_5_6_5,
  output        io_maskOut_5_6_6,
  output        io_maskOut_5_6_7,
  output        io_maskOut_5_7_0,
  output        io_maskOut_5_7_1,
  output        io_maskOut_5_7_2,
  output        io_maskOut_5_7_3,
  output        io_maskOut_5_7_4,
  output        io_maskOut_5_7_5,
  output        io_maskOut_5_7_6,
  output        io_maskOut_5_7_7,
  output        io_maskOut_6_0_0,
  output        io_maskOut_6_0_1,
  output        io_maskOut_6_0_2,
  output        io_maskOut_6_0_3,
  output        io_maskOut_6_0_4,
  output        io_maskOut_6_0_5,
  output        io_maskOut_6_0_6,
  output        io_maskOut_6_0_7,
  output        io_maskOut_6_1_0,
  output        io_maskOut_6_1_1,
  output        io_maskOut_6_1_2,
  output        io_maskOut_6_1_3,
  output        io_maskOut_6_1_4,
  output        io_maskOut_6_1_5,
  output        io_maskOut_6_1_6,
  output        io_maskOut_6_1_7,
  output        io_maskOut_6_2_0,
  output        io_maskOut_6_2_1,
  output        io_maskOut_6_2_2,
  output        io_maskOut_6_2_3,
  output        io_maskOut_6_2_4,
  output        io_maskOut_6_2_5,
  output        io_maskOut_6_2_6,
  output        io_maskOut_6_2_7,
  output        io_maskOut_6_3_0,
  output        io_maskOut_6_3_1,
  output        io_maskOut_6_3_2,
  output        io_maskOut_6_3_3,
  output        io_maskOut_6_3_4,
  output        io_maskOut_6_3_5,
  output        io_maskOut_6_3_6,
  output        io_maskOut_6_3_7,
  output        io_maskOut_6_4_0,
  output        io_maskOut_6_4_1,
  output        io_maskOut_6_4_2,
  output        io_maskOut_6_4_3,
  output        io_maskOut_6_4_4,
  output        io_maskOut_6_4_5,
  output        io_maskOut_6_4_6,
  output        io_maskOut_6_4_7,
  output        io_maskOut_6_5_0,
  output        io_maskOut_6_5_1,
  output        io_maskOut_6_5_2,
  output        io_maskOut_6_5_3,
  output        io_maskOut_6_5_4,
  output        io_maskOut_6_5_5,
  output        io_maskOut_6_5_6,
  output        io_maskOut_6_5_7,
  output        io_maskOut_6_6_0,
  output        io_maskOut_6_6_1,
  output        io_maskOut_6_6_2,
  output        io_maskOut_6_6_3,
  output        io_maskOut_6_6_4,
  output        io_maskOut_6_6_5,
  output        io_maskOut_6_6_6,
  output        io_maskOut_6_6_7,
  output        io_maskOut_6_7_0,
  output        io_maskOut_6_7_1,
  output        io_maskOut_6_7_2,
  output        io_maskOut_6_7_3,
  output        io_maskOut_6_7_4,
  output        io_maskOut_6_7_5,
  output        io_maskOut_6_7_6,
  output        io_maskOut_6_7_7,
  output        io_maskOut_7_0_0,
  output        io_maskOut_7_0_1,
  output        io_maskOut_7_0_2,
  output        io_maskOut_7_0_3,
  output        io_maskOut_7_0_4,
  output        io_maskOut_7_0_5,
  output        io_maskOut_7_0_6,
  output        io_maskOut_7_0_7,
  output        io_maskOut_7_1_0,
  output        io_maskOut_7_1_1,
  output        io_maskOut_7_1_2,
  output        io_maskOut_7_1_3,
  output        io_maskOut_7_1_4,
  output        io_maskOut_7_1_5,
  output        io_maskOut_7_1_6,
  output        io_maskOut_7_1_7,
  output        io_maskOut_7_2_0,
  output        io_maskOut_7_2_1,
  output        io_maskOut_7_2_2,
  output        io_maskOut_7_2_3,
  output        io_maskOut_7_2_4,
  output        io_maskOut_7_2_5,
  output        io_maskOut_7_2_6,
  output        io_maskOut_7_2_7,
  output        io_maskOut_7_3_0,
  output        io_maskOut_7_3_1,
  output        io_maskOut_7_3_2,
  output        io_maskOut_7_3_3,
  output        io_maskOut_7_3_4,
  output        io_maskOut_7_3_5,
  output        io_maskOut_7_3_6,
  output        io_maskOut_7_3_7,
  output        io_maskOut_7_4_0,
  output        io_maskOut_7_4_1,
  output        io_maskOut_7_4_2,
  output        io_maskOut_7_4_3,
  output        io_maskOut_7_4_4,
  output        io_maskOut_7_4_5,
  output        io_maskOut_7_4_6,
  output        io_maskOut_7_4_7,
  output        io_maskOut_7_5_0,
  output        io_maskOut_7_5_1,
  output        io_maskOut_7_5_2,
  output        io_maskOut_7_5_3,
  output        io_maskOut_7_5_4,
  output        io_maskOut_7_5_5,
  output        io_maskOut_7_5_6,
  output        io_maskOut_7_5_7,
  output        io_maskOut_7_6_0,
  output        io_maskOut_7_6_1,
  output        io_maskOut_7_6_2,
  output        io_maskOut_7_6_3,
  output        io_maskOut_7_6_4,
  output        io_maskOut_7_6_5,
  output        io_maskOut_7_6_6,
  output        io_maskOut_7_6_7,
  output        io_maskOut_7_7_0,
  output        io_maskOut_7_7_1,
  output        io_maskOut_7_7_2,
  output        io_maskOut_7_7_3,
  output        io_maskOut_7_7_4,
  output        io_maskOut_7_7_5,
  output        io_maskOut_7_7_6,
  output        io_maskOut_7_7_7,
  output        io_maskOut_8_0_0,
  output        io_maskOut_8_0_1,
  output        io_maskOut_8_0_2,
  output        io_maskOut_8_0_3,
  output        io_maskOut_8_0_4,
  output        io_maskOut_8_0_5,
  output        io_maskOut_8_0_6,
  output        io_maskOut_8_0_7,
  output        io_maskOut_8_1_0,
  output        io_maskOut_8_1_1,
  output        io_maskOut_8_1_2,
  output        io_maskOut_8_1_3,
  output        io_maskOut_8_1_4,
  output        io_maskOut_8_1_5,
  output        io_maskOut_8_1_6,
  output        io_maskOut_8_1_7,
  output        io_maskOut_8_2_0,
  output        io_maskOut_8_2_1,
  output        io_maskOut_8_2_2,
  output        io_maskOut_8_2_3,
  output        io_maskOut_8_2_4,
  output        io_maskOut_8_2_5,
  output        io_maskOut_8_2_6,
  output        io_maskOut_8_2_7,
  output        io_maskOut_8_3_0,
  output        io_maskOut_8_3_1,
  output        io_maskOut_8_3_2,
  output        io_maskOut_8_3_3,
  output        io_maskOut_8_3_4,
  output        io_maskOut_8_3_5,
  output        io_maskOut_8_3_6,
  output        io_maskOut_8_3_7,
  output        io_maskOut_8_4_0,
  output        io_maskOut_8_4_1,
  output        io_maskOut_8_4_2,
  output        io_maskOut_8_4_3,
  output        io_maskOut_8_4_4,
  output        io_maskOut_8_4_5,
  output        io_maskOut_8_4_6,
  output        io_maskOut_8_4_7,
  output        io_maskOut_8_5_0,
  output        io_maskOut_8_5_1,
  output        io_maskOut_8_5_2,
  output        io_maskOut_8_5_3,
  output        io_maskOut_8_5_4,
  output        io_maskOut_8_5_5,
  output        io_maskOut_8_5_6,
  output        io_maskOut_8_5_7,
  output        io_maskOut_8_6_0,
  output        io_maskOut_8_6_1,
  output        io_maskOut_8_6_2,
  output        io_maskOut_8_6_3,
  output        io_maskOut_8_6_4,
  output        io_maskOut_8_6_5,
  output        io_maskOut_8_6_6,
  output        io_maskOut_8_6_7,
  output        io_maskOut_8_7_0,
  output        io_maskOut_8_7_1,
  output        io_maskOut_8_7_2,
  output        io_maskOut_8_7_3,
  output        io_maskOut_8_7_4,
  output        io_maskOut_8_7_5,
  output        io_maskOut_8_7_6,
  output        io_maskOut_8_7_7,
  output        io_maskOut_9_0_0,
  output        io_maskOut_9_0_1,
  output        io_maskOut_9_0_2,
  output        io_maskOut_9_0_3,
  output        io_maskOut_9_0_4,
  output        io_maskOut_9_0_5,
  output        io_maskOut_9_0_6,
  output        io_maskOut_9_0_7,
  output        io_maskOut_9_1_0,
  output        io_maskOut_9_1_1,
  output        io_maskOut_9_1_2,
  output        io_maskOut_9_1_3,
  output        io_maskOut_9_1_4,
  output        io_maskOut_9_1_5,
  output        io_maskOut_9_1_6,
  output        io_maskOut_9_1_7,
  output        io_maskOut_9_2_0,
  output        io_maskOut_9_2_1,
  output        io_maskOut_9_2_2,
  output        io_maskOut_9_2_3,
  output        io_maskOut_9_2_4,
  output        io_maskOut_9_2_5,
  output        io_maskOut_9_2_6,
  output        io_maskOut_9_2_7,
  output        io_maskOut_9_3_0,
  output        io_maskOut_9_3_1,
  output        io_maskOut_9_3_2,
  output        io_maskOut_9_3_3,
  output        io_maskOut_9_3_4,
  output        io_maskOut_9_3_5,
  output        io_maskOut_9_3_6,
  output        io_maskOut_9_3_7,
  output        io_maskOut_9_4_0,
  output        io_maskOut_9_4_1,
  output        io_maskOut_9_4_2,
  output        io_maskOut_9_4_3,
  output        io_maskOut_9_4_4,
  output        io_maskOut_9_4_5,
  output        io_maskOut_9_4_6,
  output        io_maskOut_9_4_7,
  output        io_maskOut_9_5_0,
  output        io_maskOut_9_5_1,
  output        io_maskOut_9_5_2,
  output        io_maskOut_9_5_3,
  output        io_maskOut_9_5_4,
  output        io_maskOut_9_5_5,
  output        io_maskOut_9_5_6,
  output        io_maskOut_9_5_7,
  output        io_maskOut_9_6_0,
  output        io_maskOut_9_6_1,
  output        io_maskOut_9_6_2,
  output        io_maskOut_9_6_3,
  output        io_maskOut_9_6_4,
  output        io_maskOut_9_6_5,
  output        io_maskOut_9_6_6,
  output        io_maskOut_9_6_7,
  output        io_maskOut_9_7_0,
  output        io_maskOut_9_7_1,
  output        io_maskOut_9_7_2,
  output        io_maskOut_9_7_3,
  output        io_maskOut_9_7_4,
  output        io_maskOut_9_7_5,
  output        io_maskOut_9_7_6,
  output        io_maskOut_9_7_7,
  output        io_maskOut_10_0_0,
  output        io_maskOut_10_0_1,
  output        io_maskOut_10_0_2,
  output        io_maskOut_10_0_3,
  output        io_maskOut_10_0_4,
  output        io_maskOut_10_0_5,
  output        io_maskOut_10_0_6,
  output        io_maskOut_10_0_7,
  output        io_maskOut_10_1_0,
  output        io_maskOut_10_1_1,
  output        io_maskOut_10_1_2,
  output        io_maskOut_10_1_3,
  output        io_maskOut_10_1_4,
  output        io_maskOut_10_1_5,
  output        io_maskOut_10_1_6,
  output        io_maskOut_10_1_7,
  output        io_maskOut_10_2_0,
  output        io_maskOut_10_2_1,
  output        io_maskOut_10_2_2,
  output        io_maskOut_10_2_3,
  output        io_maskOut_10_2_4,
  output        io_maskOut_10_2_5,
  output        io_maskOut_10_2_6,
  output        io_maskOut_10_2_7,
  output        io_maskOut_10_3_0,
  output        io_maskOut_10_3_1,
  output        io_maskOut_10_3_2,
  output        io_maskOut_10_3_3,
  output        io_maskOut_10_3_4,
  output        io_maskOut_10_3_5,
  output        io_maskOut_10_3_6,
  output        io_maskOut_10_3_7,
  output        io_maskOut_10_4_0,
  output        io_maskOut_10_4_1,
  output        io_maskOut_10_4_2,
  output        io_maskOut_10_4_3,
  output        io_maskOut_10_4_4,
  output        io_maskOut_10_4_5,
  output        io_maskOut_10_4_6,
  output        io_maskOut_10_4_7,
  output        io_maskOut_10_5_0,
  output        io_maskOut_10_5_1,
  output        io_maskOut_10_5_2,
  output        io_maskOut_10_5_3,
  output        io_maskOut_10_5_4,
  output        io_maskOut_10_5_5,
  output        io_maskOut_10_5_6,
  output        io_maskOut_10_5_7,
  output        io_maskOut_10_6_0,
  output        io_maskOut_10_6_1,
  output        io_maskOut_10_6_2,
  output        io_maskOut_10_6_3,
  output        io_maskOut_10_6_4,
  output        io_maskOut_10_6_5,
  output        io_maskOut_10_6_6,
  output        io_maskOut_10_6_7,
  output        io_maskOut_10_7_0,
  output        io_maskOut_10_7_1,
  output        io_maskOut_10_7_2,
  output        io_maskOut_10_7_3,
  output        io_maskOut_10_7_4,
  output        io_maskOut_10_7_5,
  output        io_maskOut_10_7_6,
  output        io_maskOut_10_7_7,
  output        io_maskOut_11_0_0,
  output        io_maskOut_11_0_1,
  output        io_maskOut_11_0_2,
  output        io_maskOut_11_0_3,
  output        io_maskOut_11_0_4,
  output        io_maskOut_11_0_5,
  output        io_maskOut_11_0_6,
  output        io_maskOut_11_0_7,
  output        io_maskOut_11_1_0,
  output        io_maskOut_11_1_1,
  output        io_maskOut_11_1_2,
  output        io_maskOut_11_1_3,
  output        io_maskOut_11_1_4,
  output        io_maskOut_11_1_5,
  output        io_maskOut_11_1_6,
  output        io_maskOut_11_1_7,
  output        io_maskOut_11_2_0,
  output        io_maskOut_11_2_1,
  output        io_maskOut_11_2_2,
  output        io_maskOut_11_2_3,
  output        io_maskOut_11_2_4,
  output        io_maskOut_11_2_5,
  output        io_maskOut_11_2_6,
  output        io_maskOut_11_2_7,
  output        io_maskOut_11_3_0,
  output        io_maskOut_11_3_1,
  output        io_maskOut_11_3_2,
  output        io_maskOut_11_3_3,
  output        io_maskOut_11_3_4,
  output        io_maskOut_11_3_5,
  output        io_maskOut_11_3_6,
  output        io_maskOut_11_3_7,
  output        io_maskOut_11_4_0,
  output        io_maskOut_11_4_1,
  output        io_maskOut_11_4_2,
  output        io_maskOut_11_4_3,
  output        io_maskOut_11_4_4,
  output        io_maskOut_11_4_5,
  output        io_maskOut_11_4_6,
  output        io_maskOut_11_4_7,
  output        io_maskOut_11_5_0,
  output        io_maskOut_11_5_1,
  output        io_maskOut_11_5_2,
  output        io_maskOut_11_5_3,
  output        io_maskOut_11_5_4,
  output        io_maskOut_11_5_5,
  output        io_maskOut_11_5_6,
  output        io_maskOut_11_5_7,
  output        io_maskOut_11_6_0,
  output        io_maskOut_11_6_1,
  output        io_maskOut_11_6_2,
  output        io_maskOut_11_6_3,
  output        io_maskOut_11_6_4,
  output        io_maskOut_11_6_5,
  output        io_maskOut_11_6_6,
  output        io_maskOut_11_6_7,
  output        io_maskOut_11_7_0,
  output        io_maskOut_11_7_1,
  output        io_maskOut_11_7_2,
  output        io_maskOut_11_7_3,
  output        io_maskOut_11_7_4,
  output        io_maskOut_11_7_5,
  output        io_maskOut_11_7_6,
  output        io_maskOut_11_7_7,
  output        io_maskOut_12_0_0,
  output        io_maskOut_12_0_1,
  output        io_maskOut_12_0_2,
  output        io_maskOut_12_0_3,
  output        io_maskOut_12_0_4,
  output        io_maskOut_12_0_5,
  output        io_maskOut_12_0_6,
  output        io_maskOut_12_0_7,
  output        io_maskOut_12_1_0,
  output        io_maskOut_12_1_1,
  output        io_maskOut_12_1_2,
  output        io_maskOut_12_1_3,
  output        io_maskOut_12_1_4,
  output        io_maskOut_12_1_5,
  output        io_maskOut_12_1_6,
  output        io_maskOut_12_1_7,
  output        io_maskOut_12_2_0,
  output        io_maskOut_12_2_1,
  output        io_maskOut_12_2_2,
  output        io_maskOut_12_2_3,
  output        io_maskOut_12_2_4,
  output        io_maskOut_12_2_5,
  output        io_maskOut_12_2_6,
  output        io_maskOut_12_2_7,
  output        io_maskOut_12_3_0,
  output        io_maskOut_12_3_1,
  output        io_maskOut_12_3_2,
  output        io_maskOut_12_3_3,
  output        io_maskOut_12_3_4,
  output        io_maskOut_12_3_5,
  output        io_maskOut_12_3_6,
  output        io_maskOut_12_3_7,
  output        io_maskOut_12_4_0,
  output        io_maskOut_12_4_1,
  output        io_maskOut_12_4_2,
  output        io_maskOut_12_4_3,
  output        io_maskOut_12_4_4,
  output        io_maskOut_12_4_5,
  output        io_maskOut_12_4_6,
  output        io_maskOut_12_4_7,
  output        io_maskOut_12_5_0,
  output        io_maskOut_12_5_1,
  output        io_maskOut_12_5_2,
  output        io_maskOut_12_5_3,
  output        io_maskOut_12_5_4,
  output        io_maskOut_12_5_5,
  output        io_maskOut_12_5_6,
  output        io_maskOut_12_5_7,
  output        io_maskOut_12_6_0,
  output        io_maskOut_12_6_1,
  output        io_maskOut_12_6_2,
  output        io_maskOut_12_6_3,
  output        io_maskOut_12_6_4,
  output        io_maskOut_12_6_5,
  output        io_maskOut_12_6_6,
  output        io_maskOut_12_6_7,
  output        io_maskOut_12_7_0,
  output        io_maskOut_12_7_1,
  output        io_maskOut_12_7_2,
  output        io_maskOut_12_7_3,
  output        io_maskOut_12_7_4,
  output        io_maskOut_12_7_5,
  output        io_maskOut_12_7_6,
  output        io_maskOut_12_7_7,
  output        io_maskOut_13_0_0,
  output        io_maskOut_13_0_1,
  output        io_maskOut_13_0_2,
  output        io_maskOut_13_0_3,
  output        io_maskOut_13_0_4,
  output        io_maskOut_13_0_5,
  output        io_maskOut_13_0_6,
  output        io_maskOut_13_0_7,
  output        io_maskOut_13_1_0,
  output        io_maskOut_13_1_1,
  output        io_maskOut_13_1_2,
  output        io_maskOut_13_1_3,
  output        io_maskOut_13_1_4,
  output        io_maskOut_13_1_5,
  output        io_maskOut_13_1_6,
  output        io_maskOut_13_1_7,
  output        io_maskOut_13_2_0,
  output        io_maskOut_13_2_1,
  output        io_maskOut_13_2_2,
  output        io_maskOut_13_2_3,
  output        io_maskOut_13_2_4,
  output        io_maskOut_13_2_5,
  output        io_maskOut_13_2_6,
  output        io_maskOut_13_2_7,
  output        io_maskOut_13_3_0,
  output        io_maskOut_13_3_1,
  output        io_maskOut_13_3_2,
  output        io_maskOut_13_3_3,
  output        io_maskOut_13_3_4,
  output        io_maskOut_13_3_5,
  output        io_maskOut_13_3_6,
  output        io_maskOut_13_3_7,
  output        io_maskOut_13_4_0,
  output        io_maskOut_13_4_1,
  output        io_maskOut_13_4_2,
  output        io_maskOut_13_4_3,
  output        io_maskOut_13_4_4,
  output        io_maskOut_13_4_5,
  output        io_maskOut_13_4_6,
  output        io_maskOut_13_4_7,
  output        io_maskOut_13_5_0,
  output        io_maskOut_13_5_1,
  output        io_maskOut_13_5_2,
  output        io_maskOut_13_5_3,
  output        io_maskOut_13_5_4,
  output        io_maskOut_13_5_5,
  output        io_maskOut_13_5_6,
  output        io_maskOut_13_5_7,
  output        io_maskOut_13_6_0,
  output        io_maskOut_13_6_1,
  output        io_maskOut_13_6_2,
  output        io_maskOut_13_6_3,
  output        io_maskOut_13_6_4,
  output        io_maskOut_13_6_5,
  output        io_maskOut_13_6_6,
  output        io_maskOut_13_6_7,
  output        io_maskOut_13_7_0,
  output        io_maskOut_13_7_1,
  output        io_maskOut_13_7_2,
  output        io_maskOut_13_7_3,
  output        io_maskOut_13_7_4,
  output        io_maskOut_13_7_5,
  output        io_maskOut_13_7_6,
  output        io_maskOut_13_7_7,
  output        io_maskOut_14_0_0,
  output        io_maskOut_14_0_1,
  output        io_maskOut_14_0_2,
  output        io_maskOut_14_0_3,
  output        io_maskOut_14_0_4,
  output        io_maskOut_14_0_5,
  output        io_maskOut_14_0_6,
  output        io_maskOut_14_0_7,
  output        io_maskOut_14_1_0,
  output        io_maskOut_14_1_1,
  output        io_maskOut_14_1_2,
  output        io_maskOut_14_1_3,
  output        io_maskOut_14_1_4,
  output        io_maskOut_14_1_5,
  output        io_maskOut_14_1_6,
  output        io_maskOut_14_1_7,
  output        io_maskOut_14_2_0,
  output        io_maskOut_14_2_1,
  output        io_maskOut_14_2_2,
  output        io_maskOut_14_2_3,
  output        io_maskOut_14_2_4,
  output        io_maskOut_14_2_5,
  output        io_maskOut_14_2_6,
  output        io_maskOut_14_2_7,
  output        io_maskOut_14_3_0,
  output        io_maskOut_14_3_1,
  output        io_maskOut_14_3_2,
  output        io_maskOut_14_3_3,
  output        io_maskOut_14_3_4,
  output        io_maskOut_14_3_5,
  output        io_maskOut_14_3_6,
  output        io_maskOut_14_3_7,
  output        io_maskOut_14_4_0,
  output        io_maskOut_14_4_1,
  output        io_maskOut_14_4_2,
  output        io_maskOut_14_4_3,
  output        io_maskOut_14_4_4,
  output        io_maskOut_14_4_5,
  output        io_maskOut_14_4_6,
  output        io_maskOut_14_4_7,
  output        io_maskOut_14_5_0,
  output        io_maskOut_14_5_1,
  output        io_maskOut_14_5_2,
  output        io_maskOut_14_5_3,
  output        io_maskOut_14_5_4,
  output        io_maskOut_14_5_5,
  output        io_maskOut_14_5_6,
  output        io_maskOut_14_5_7,
  output        io_maskOut_14_6_0,
  output        io_maskOut_14_6_1,
  output        io_maskOut_14_6_2,
  output        io_maskOut_14_6_3,
  output        io_maskOut_14_6_4,
  output        io_maskOut_14_6_5,
  output        io_maskOut_14_6_6,
  output        io_maskOut_14_6_7,
  output        io_maskOut_14_7_0,
  output        io_maskOut_14_7_1,
  output        io_maskOut_14_7_2,
  output        io_maskOut_14_7_3,
  output        io_maskOut_14_7_4,
  output        io_maskOut_14_7_5,
  output        io_maskOut_14_7_6,
  output        io_maskOut_14_7_7,
  output        io_maskOut_15_0_0,
  output        io_maskOut_15_0_1,
  output        io_maskOut_15_0_2,
  output        io_maskOut_15_0_3,
  output        io_maskOut_15_0_4,
  output        io_maskOut_15_0_5,
  output        io_maskOut_15_0_6,
  output        io_maskOut_15_0_7,
  output        io_maskOut_15_1_0,
  output        io_maskOut_15_1_1,
  output        io_maskOut_15_1_2,
  output        io_maskOut_15_1_3,
  output        io_maskOut_15_1_4,
  output        io_maskOut_15_1_5,
  output        io_maskOut_15_1_6,
  output        io_maskOut_15_1_7,
  output        io_maskOut_15_2_0,
  output        io_maskOut_15_2_1,
  output        io_maskOut_15_2_2,
  output        io_maskOut_15_2_3,
  output        io_maskOut_15_2_4,
  output        io_maskOut_15_2_5,
  output        io_maskOut_15_2_6,
  output        io_maskOut_15_2_7,
  output        io_maskOut_15_3_0,
  output        io_maskOut_15_3_1,
  output        io_maskOut_15_3_2,
  output        io_maskOut_15_3_3,
  output        io_maskOut_15_3_4,
  output        io_maskOut_15_3_5,
  output        io_maskOut_15_3_6,
  output        io_maskOut_15_3_7,
  output        io_maskOut_15_4_0,
  output        io_maskOut_15_4_1,
  output        io_maskOut_15_4_2,
  output        io_maskOut_15_4_3,
  output        io_maskOut_15_4_4,
  output        io_maskOut_15_4_5,
  output        io_maskOut_15_4_6,
  output        io_maskOut_15_4_7,
  output        io_maskOut_15_5_0,
  output        io_maskOut_15_5_1,
  output        io_maskOut_15_5_2,
  output        io_maskOut_15_5_3,
  output        io_maskOut_15_5_4,
  output        io_maskOut_15_5_5,
  output        io_maskOut_15_5_6,
  output        io_maskOut_15_5_7,
  output        io_maskOut_15_6_0,
  output        io_maskOut_15_6_1,
  output        io_maskOut_15_6_2,
  output        io_maskOut_15_6_3,
  output        io_maskOut_15_6_4,
  output        io_maskOut_15_6_5,
  output        io_maskOut_15_6_6,
  output        io_maskOut_15_6_7,
  output        io_maskOut_15_7_0,
  output        io_maskOut_15_7_1,
  output        io_maskOut_15_7_2,
  output        io_maskOut_15_7_3,
  output        io_maskOut_15_7_4,
  output        io_maskOut_15_7_5,
  output        io_maskOut_15_7_6,
  output        io_maskOut_15_7_7
);
  reg [7:0] data_0_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_0_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_1_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_2_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_3_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_4_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_5_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_6_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_7_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_8_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_9_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_10_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_11_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_12_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_13_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_14_7_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_0_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_1_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_2_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_3_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_4_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_5_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_6_7; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_0; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_1; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_2; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_3; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_4; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_5; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_6; // @[Sbuffer.scala 96:17]
  reg [7:0] data_15_7_7; // @[Sbuffer.scala 96:17]
  reg  mask_0_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_0_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_1_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_2_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_3_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_4_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_5_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_6_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_7_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_8_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_9_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_10_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_11_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_12_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_13_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_14_7_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_0_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_1_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_2_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_3_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_4_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_5_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_6_7; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_0; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_1; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_2; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_3; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_4; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_5; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_6; // @[Sbuffer.scala 98:21]
  reg  mask_15_7_7; // @[Sbuffer.scala 98:21]
  reg  line_mask_clean_valid_0; // @[Sbuffer.scala 121:63]
  reg  line_mask_clean_valid_1; // @[Sbuffer.scala 121:63]
  wire [7:0] line_mask_clean_line_hi = io_maskFlushReq_0_bits_wvec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] line_mask_clean_line_lo = io_maskFlushReq_0_bits_wvec[7:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T = |line_mask_clean_line_hi; // @[OneHot.scala 32:14]
  wire [7:0] _line_mask_clean_line_T_1 = line_mask_clean_line_hi | line_mask_clean_line_lo; // @[OneHot.scala 32:28]
  wire [3:0] line_mask_clean_line_hi_1 = _line_mask_clean_line_T_1[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] line_mask_clean_line_lo_1 = _line_mask_clean_line_T_1[3:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T_2 = |line_mask_clean_line_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _line_mask_clean_line_T_3 = line_mask_clean_line_hi_1 | line_mask_clean_line_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] line_mask_clean_line_hi_2 = _line_mask_clean_line_T_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] line_mask_clean_line_lo_2 = _line_mask_clean_line_T_3[1:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T_4 = |line_mask_clean_line_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _line_mask_clean_line_T_5 = line_mask_clean_line_hi_2 | line_mask_clean_line_lo_2; // @[OneHot.scala 32:28]
  wire [2:0] _line_mask_clean_line_T_8 = {_line_mask_clean_line_T_2,_line_mask_clean_line_T_4,_line_mask_clean_line_T_5[
    1]}; // @[Cat.scala 33:92]
  reg [3:0] line_mask_clean_line_0; // @[Sbuffer.scala 122:62]
  wire [7:0] line_mask_clean_line_hi_3 = io_maskFlushReq_1_bits_wvec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] line_mask_clean_line_lo_3 = io_maskFlushReq_1_bits_wvec[7:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T_10 = |line_mask_clean_line_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _line_mask_clean_line_T_11 = line_mask_clean_line_hi_3 | line_mask_clean_line_lo_3; // @[OneHot.scala 32:28]
  wire [3:0] line_mask_clean_line_hi_4 = _line_mask_clean_line_T_11[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] line_mask_clean_line_lo_4 = _line_mask_clean_line_T_11[3:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T_12 = |line_mask_clean_line_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _line_mask_clean_line_T_13 = line_mask_clean_line_hi_4 | line_mask_clean_line_lo_4; // @[OneHot.scala 32:28]
  wire [1:0] line_mask_clean_line_hi_5 = _line_mask_clean_line_T_13[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] line_mask_clean_line_lo_5 = _line_mask_clean_line_T_13[1:0]; // @[OneHot.scala 31:18]
  wire  _line_mask_clean_line_T_14 = |line_mask_clean_line_hi_5; // @[OneHot.scala 32:14]
  wire [1:0] _line_mask_clean_line_T_15 = line_mask_clean_line_hi_5 | line_mask_clean_line_lo_5; // @[OneHot.scala 32:28]
  wire [2:0] _line_mask_clean_line_T_18 = {_line_mask_clean_line_T_12,_line_mask_clean_line_T_14,
    _line_mask_clean_line_T_15[1]}; // @[Cat.scala 33:92]
  reg [3:0] line_mask_clean_line_1; // @[Sbuffer.scala 122:62]
  wire  _GEN_0 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_2 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_3 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_4 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_5 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_6 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_7 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_8 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_9 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_10 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_11 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_12 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_13 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_14 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_15 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_16 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_17 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_18 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_19 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_20 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_21 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_22 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_23 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_24 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_25 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_26 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_27 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_28 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_29 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_30 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_31 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_32 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_33 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_34 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_35 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_36 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_37 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_38 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_39 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_40 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_41 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_42 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_43 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_44 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_45 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_46 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_47 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_48 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_49 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_50 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_51 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_52 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_53 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_54 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_55 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_56 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_57 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_58 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_59 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_60 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_61 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_62 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_63 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_64 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_65 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_66 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_67 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_68 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_69 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_70 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_71 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_72 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_73 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_74 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_75 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_76 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_77 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_78 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_79 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_80 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_81 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_82 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_83 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_84 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_85 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_86 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_87 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_88 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_89 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_90 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_91 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_92 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_93 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_94 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_95 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_96 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_97 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_98 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_99 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_100 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_101 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_102 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_103 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_104 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_105 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_106 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_107 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_108 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_109 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_110 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_111 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_112 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_113 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_114 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_115 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_116 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_117 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_118 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_119 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_120 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_121 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_122 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_123 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_124 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_125 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_126 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_127 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_0_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_128 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_129 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_130 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_131 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_132 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_133 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_134 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_135 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_136 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_137 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_138 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_139 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_140 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_141 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_142 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_143 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_144 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_145 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_146 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_147 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_148 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_149 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_150 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_151 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_152 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_153 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_154 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_155 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_156 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_157 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_158 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_159 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_160 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_161 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_162 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_163 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_164 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_165 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_166 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_167 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_168 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_169 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_170 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_171 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_172 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_173 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_174 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_175 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_176 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_177 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_178 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_179 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_180 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_181 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_182 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_183 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_184 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_185 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_186 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_187 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_188 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_189 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_190 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_191 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_192 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_193 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_194 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_195 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_196 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_197 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_198 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_199 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_200 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_201 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_202 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_203 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_204 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_205 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_206 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_207 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_208 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_209 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_210 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_211 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_212 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_213 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_214 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_215 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_216 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_217 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_218 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_219 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_220 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_221 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_222 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_223 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_224 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_225 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_226 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_227 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_228 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_229 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_230 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_231 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_232 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_233 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_234 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_235 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_236 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_237 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_238 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_239 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_240 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_241 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_242 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_243 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_244 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_245 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_246 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_247 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_248 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_249 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_250 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_251 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_252 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_253 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_254 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_255 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_1_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_256 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_257 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_258 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_259 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_260 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_261 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_262 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_263 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_264 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_265 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_266 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_267 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_268 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_269 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_270 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_271 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_272 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_273 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_274 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_275 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_276 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_277 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_278 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_279 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_280 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_281 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_282 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_283 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_284 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_285 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_286 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_287 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_288 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_289 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_290 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_291 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_292 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_293 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_294 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_295 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_296 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_297 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_298 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_299 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_300 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_301 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_302 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_303 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_304 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_305 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_306 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_307 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_308 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_309 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_310 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_311 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_312 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_313 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_314 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_315 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_316 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_317 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_318 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_319 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_320 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_321 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_322 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_323 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_324 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_325 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_326 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_327 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_328 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_329 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_330 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_331 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_332 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_333 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_334 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_335 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_336 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_337 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_338 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_339 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_340 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_341 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_342 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_343 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_344 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_345 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_346 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_347 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_348 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_349 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_350 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_351 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_352 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_353 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_354 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_355 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_356 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_357 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_358 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_359 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_360 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_361 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_362 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_363 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_364 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_365 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_366 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_367 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_368 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_369 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_370 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_371 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_372 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_373 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_374 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_375 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_376 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_377 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_378 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_379 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_380 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_381 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_382 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_383 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_2_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_384 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_385 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_386 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_387 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_388 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_389 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_390 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_391 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_392 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_393 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_394 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_395 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_396 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_397 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_398 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_399 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_400 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_401 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_402 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_403 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_404 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_405 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_406 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_407 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_408 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_409 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_410 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_411 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_412 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_413 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_414 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_415 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_416 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_417 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_418 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_419 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_420 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_421 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_422 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_423 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_424 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_425 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_426 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_427 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_428 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_429 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_430 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_431 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_432 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_433 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_434 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_435 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_436 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_437 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_438 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_439 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_440 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_441 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_442 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_443 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_444 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_445 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_446 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_447 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_448 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_449 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_450 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_451 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_452 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_453 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_454 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_455 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_456 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_457 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_458 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_459 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_460 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_461 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_462 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_463 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_464 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_465 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_466 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_467 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_468 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_469 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_470 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_471 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_472 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_473 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_474 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_475 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_476 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_477 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_478 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_479 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_480 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_481 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_482 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_483 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_484 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_485 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_486 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_487 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_488 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_489 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_490 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_491 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_492 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_493 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_494 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_495 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_496 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_497 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_498 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_499 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_500 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_501 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_502 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_503 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_504 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_505 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_506 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_507 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_508 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_509 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_510 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_511 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_3_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_512 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_513 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_514 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_515 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_516 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_517 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_518 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_519 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_520 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_521 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_522 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_523 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_524 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_525 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_526 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_527 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_528 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_529 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_530 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_531 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_532 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_533 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_534 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_535 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_536 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_537 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_538 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_539 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_540 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_541 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_542 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_543 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_544 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_545 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_546 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_547 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_548 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_549 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_550 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_551 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_552 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_553 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_554 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_555 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_556 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_557 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_558 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_559 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_560 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_561 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_562 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_563 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_564 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_565 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_566 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_567 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_568 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_569 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_570 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_571 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_572 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_573 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_574 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_575 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_576 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_577 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_578 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_579 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_580 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_581 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_582 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_583 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_584 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_585 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_586 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_587 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_588 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_589 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_590 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_591 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_592 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_593 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_594 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_595 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_596 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_597 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_598 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_599 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_600 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_601 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_602 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_603 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_604 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_605 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_606 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_607 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_608 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_609 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_610 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_611 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_612 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_613 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_614 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_615 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_616 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_617 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_618 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_619 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_620 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_621 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_622 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_623 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_624 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_625 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_626 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_627 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_628 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_629 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_630 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_631 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_632 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_633 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_634 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_635 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_636 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_637 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_638 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_639 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_4_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_640 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_641 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_642 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_643 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_644 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_645 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_646 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_647 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_648 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_649 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_650 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_651 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_652 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_653 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_654 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_655 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_656 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_657 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_658 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_659 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_660 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_661 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_662 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_663 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_664 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_665 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_666 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_667 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_668 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_669 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_670 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_671 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_672 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_673 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_674 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_675 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_676 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_677 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_678 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_679 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_680 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_681 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_682 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_683 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_684 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_685 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_686 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_687 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_688 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_689 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_690 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_691 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_692 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_693 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_694 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_695 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_696 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_697 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_698 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_699 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_700 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_701 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_702 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_703 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_704 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_705 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_706 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_707 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_708 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_709 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_710 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_711 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_712 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_713 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_714 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_715 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_716 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_717 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_718 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_719 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_720 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_721 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_722 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_723 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_724 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_725 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_726 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_727 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_728 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_729 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_730 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_731 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_732 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_733 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_734 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_735 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_736 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_737 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_738 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_739 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_740 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_741 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_742 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_743 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_744 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_745 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_746 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_747 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_748 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_749 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_750 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_751 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_752 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_753 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_754 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_755 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_756 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_757 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_758 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_759 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_760 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_761 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_762 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_763 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_764 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_765 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_766 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_767 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_5_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_768 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_769 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_770 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_771 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_772 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_773 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_774 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_775 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_776 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_777 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_778 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_779 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_780 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_781 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_782 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_783 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_784 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_785 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_786 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_787 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_788 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_789 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_790 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_791 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_792 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_793 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_794 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_795 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_796 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_797 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_798 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_799 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_800 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_801 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_802 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_803 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_804 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_805 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_806 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_807 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_808 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_809 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_810 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_811 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_812 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_813 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_814 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_815 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_816 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_817 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_818 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_819 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_820 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_821 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_822 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_823 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_824 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_825 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_826 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_827 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_828 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_829 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_830 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_831 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_832 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_833 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_834 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_835 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_836 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_837 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_838 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_839 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_840 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_841 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_842 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_843 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_844 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_845 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_846 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_847 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_848 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_849 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_850 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_851 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_852 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_853 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_854 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_855 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_856 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_857 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_858 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_859 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_860 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_861 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_862 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_863 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_864 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_865 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_866 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_867 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_868 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_869 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_870 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_871 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_872 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_873 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_874 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_875 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_876 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_877 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_878 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_879 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_880 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_881 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_882 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_883 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_884 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_885 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_886 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_887 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_888 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_889 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_890 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_891 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_892 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_893 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_894 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_895 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_6_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_896 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_897 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_898 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_899 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_900 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_901 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_902 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_903 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_904 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_905 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_906 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_907 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_908 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_909 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_910 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_911 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_0; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_912 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_913 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_914 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_915 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_916 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_917 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_918 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_919 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_920 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_921 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_922 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_923 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_924 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_925 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_926 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_927 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_1; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_928 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_929 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_930 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_931 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_932 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_933 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_934 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_935 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_936 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_937 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_938 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_939 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_940 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_941 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_942 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_943 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_2; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_944 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_945 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_946 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_947 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_948 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_949 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_950 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_951 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_952 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_953 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_954 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_955 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_956 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_957 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_958 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_959 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_3; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_960 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_961 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_962 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_963 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_964 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_965 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_966 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_967 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_968 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_969 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_970 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_971 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_972 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_973 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_974 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_975 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_4; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_976 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_977 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_978 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_979 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_980 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_981 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_982 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_983 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_984 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_985 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_986 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_987 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_988 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_989 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_990 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_991 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_5; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_992 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_993 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_994 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_995 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_996 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_997 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_998 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_999 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1000 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1001 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1002 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1003 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1004 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1005 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1006 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1007 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_6; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1008 = 4'h0 == line_mask_clean_line_0 ? 1'h0 : mask_0_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1009 = 4'h1 == line_mask_clean_line_0 ? 1'h0 : mask_1_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1010 = 4'h2 == line_mask_clean_line_0 ? 1'h0 : mask_2_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1011 = 4'h3 == line_mask_clean_line_0 ? 1'h0 : mask_3_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1012 = 4'h4 == line_mask_clean_line_0 ? 1'h0 : mask_4_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1013 = 4'h5 == line_mask_clean_line_0 ? 1'h0 : mask_5_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1014 = 4'h6 == line_mask_clean_line_0 ? 1'h0 : mask_6_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1015 = 4'h7 == line_mask_clean_line_0 ? 1'h0 : mask_7_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1016 = 4'h8 == line_mask_clean_line_0 ? 1'h0 : mask_8_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1017 = 4'h9 == line_mask_clean_line_0 ? 1'h0 : mask_9_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1018 = 4'ha == line_mask_clean_line_0 ? 1'h0 : mask_10_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1019 = 4'hb == line_mask_clean_line_0 ? 1'h0 : mask_11_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1020 = 4'hc == line_mask_clean_line_0 ? 1'h0 : mask_12_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1021 = 4'hd == line_mask_clean_line_0 ? 1'h0 : mask_13_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1022 = 4'he == line_mask_clean_line_0 ? 1'h0 : mask_14_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1023 = 4'hf == line_mask_clean_line_0 ? 1'h0 : mask_15_7_7; // @[Sbuffer.scala 137:{34,34} 98:21]
  wire  _GEN_1024 = line_mask_clean_valid_0 ? _GEN_0 : mask_0_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1025 = line_mask_clean_valid_0 ? _GEN_1 : mask_1_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1026 = line_mask_clean_valid_0 ? _GEN_2 : mask_2_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1027 = line_mask_clean_valid_0 ? _GEN_3 : mask_3_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1028 = line_mask_clean_valid_0 ? _GEN_4 : mask_4_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1029 = line_mask_clean_valid_0 ? _GEN_5 : mask_5_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1030 = line_mask_clean_valid_0 ? _GEN_6 : mask_6_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1031 = line_mask_clean_valid_0 ? _GEN_7 : mask_7_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1032 = line_mask_clean_valid_0 ? _GEN_8 : mask_8_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1033 = line_mask_clean_valid_0 ? _GEN_9 : mask_9_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1034 = line_mask_clean_valid_0 ? _GEN_10 : mask_10_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1035 = line_mask_clean_valid_0 ? _GEN_11 : mask_11_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1036 = line_mask_clean_valid_0 ? _GEN_12 : mask_12_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1037 = line_mask_clean_valid_0 ? _GEN_13 : mask_13_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1038 = line_mask_clean_valid_0 ? _GEN_14 : mask_14_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1039 = line_mask_clean_valid_0 ? _GEN_15 : mask_15_0_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1040 = line_mask_clean_valid_0 ? _GEN_16 : mask_0_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1041 = line_mask_clean_valid_0 ? _GEN_17 : mask_1_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1042 = line_mask_clean_valid_0 ? _GEN_18 : mask_2_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1043 = line_mask_clean_valid_0 ? _GEN_19 : mask_3_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1044 = line_mask_clean_valid_0 ? _GEN_20 : mask_4_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1045 = line_mask_clean_valid_0 ? _GEN_21 : mask_5_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1046 = line_mask_clean_valid_0 ? _GEN_22 : mask_6_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1047 = line_mask_clean_valid_0 ? _GEN_23 : mask_7_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1048 = line_mask_clean_valid_0 ? _GEN_24 : mask_8_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1049 = line_mask_clean_valid_0 ? _GEN_25 : mask_9_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1050 = line_mask_clean_valid_0 ? _GEN_26 : mask_10_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1051 = line_mask_clean_valid_0 ? _GEN_27 : mask_11_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1052 = line_mask_clean_valid_0 ? _GEN_28 : mask_12_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1053 = line_mask_clean_valid_0 ? _GEN_29 : mask_13_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1054 = line_mask_clean_valid_0 ? _GEN_30 : mask_14_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1055 = line_mask_clean_valid_0 ? _GEN_31 : mask_15_0_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1056 = line_mask_clean_valid_0 ? _GEN_32 : mask_0_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1057 = line_mask_clean_valid_0 ? _GEN_33 : mask_1_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1058 = line_mask_clean_valid_0 ? _GEN_34 : mask_2_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1059 = line_mask_clean_valid_0 ? _GEN_35 : mask_3_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1060 = line_mask_clean_valid_0 ? _GEN_36 : mask_4_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1061 = line_mask_clean_valid_0 ? _GEN_37 : mask_5_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1062 = line_mask_clean_valid_0 ? _GEN_38 : mask_6_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1063 = line_mask_clean_valid_0 ? _GEN_39 : mask_7_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1064 = line_mask_clean_valid_0 ? _GEN_40 : mask_8_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1065 = line_mask_clean_valid_0 ? _GEN_41 : mask_9_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1066 = line_mask_clean_valid_0 ? _GEN_42 : mask_10_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1067 = line_mask_clean_valid_0 ? _GEN_43 : mask_11_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1068 = line_mask_clean_valid_0 ? _GEN_44 : mask_12_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1069 = line_mask_clean_valid_0 ? _GEN_45 : mask_13_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1070 = line_mask_clean_valid_0 ? _GEN_46 : mask_14_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1071 = line_mask_clean_valid_0 ? _GEN_47 : mask_15_0_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1072 = line_mask_clean_valid_0 ? _GEN_48 : mask_0_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1073 = line_mask_clean_valid_0 ? _GEN_49 : mask_1_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1074 = line_mask_clean_valid_0 ? _GEN_50 : mask_2_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1075 = line_mask_clean_valid_0 ? _GEN_51 : mask_3_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1076 = line_mask_clean_valid_0 ? _GEN_52 : mask_4_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1077 = line_mask_clean_valid_0 ? _GEN_53 : mask_5_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1078 = line_mask_clean_valid_0 ? _GEN_54 : mask_6_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1079 = line_mask_clean_valid_0 ? _GEN_55 : mask_7_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1080 = line_mask_clean_valid_0 ? _GEN_56 : mask_8_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1081 = line_mask_clean_valid_0 ? _GEN_57 : mask_9_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1082 = line_mask_clean_valid_0 ? _GEN_58 : mask_10_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1083 = line_mask_clean_valid_0 ? _GEN_59 : mask_11_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1084 = line_mask_clean_valid_0 ? _GEN_60 : mask_12_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1085 = line_mask_clean_valid_0 ? _GEN_61 : mask_13_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1086 = line_mask_clean_valid_0 ? _GEN_62 : mask_14_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1087 = line_mask_clean_valid_0 ? _GEN_63 : mask_15_0_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1088 = line_mask_clean_valid_0 ? _GEN_64 : mask_0_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1089 = line_mask_clean_valid_0 ? _GEN_65 : mask_1_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1090 = line_mask_clean_valid_0 ? _GEN_66 : mask_2_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1091 = line_mask_clean_valid_0 ? _GEN_67 : mask_3_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1092 = line_mask_clean_valid_0 ? _GEN_68 : mask_4_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1093 = line_mask_clean_valid_0 ? _GEN_69 : mask_5_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1094 = line_mask_clean_valid_0 ? _GEN_70 : mask_6_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1095 = line_mask_clean_valid_0 ? _GEN_71 : mask_7_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1096 = line_mask_clean_valid_0 ? _GEN_72 : mask_8_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1097 = line_mask_clean_valid_0 ? _GEN_73 : mask_9_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1098 = line_mask_clean_valid_0 ? _GEN_74 : mask_10_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1099 = line_mask_clean_valid_0 ? _GEN_75 : mask_11_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1100 = line_mask_clean_valid_0 ? _GEN_76 : mask_12_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1101 = line_mask_clean_valid_0 ? _GEN_77 : mask_13_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1102 = line_mask_clean_valid_0 ? _GEN_78 : mask_14_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1103 = line_mask_clean_valid_0 ? _GEN_79 : mask_15_0_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1104 = line_mask_clean_valid_0 ? _GEN_80 : mask_0_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1105 = line_mask_clean_valid_0 ? _GEN_81 : mask_1_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1106 = line_mask_clean_valid_0 ? _GEN_82 : mask_2_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1107 = line_mask_clean_valid_0 ? _GEN_83 : mask_3_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1108 = line_mask_clean_valid_0 ? _GEN_84 : mask_4_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1109 = line_mask_clean_valid_0 ? _GEN_85 : mask_5_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1110 = line_mask_clean_valid_0 ? _GEN_86 : mask_6_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1111 = line_mask_clean_valid_0 ? _GEN_87 : mask_7_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1112 = line_mask_clean_valid_0 ? _GEN_88 : mask_8_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1113 = line_mask_clean_valid_0 ? _GEN_89 : mask_9_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1114 = line_mask_clean_valid_0 ? _GEN_90 : mask_10_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1115 = line_mask_clean_valid_0 ? _GEN_91 : mask_11_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1116 = line_mask_clean_valid_0 ? _GEN_92 : mask_12_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1117 = line_mask_clean_valid_0 ? _GEN_93 : mask_13_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1118 = line_mask_clean_valid_0 ? _GEN_94 : mask_14_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1119 = line_mask_clean_valid_0 ? _GEN_95 : mask_15_0_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1120 = line_mask_clean_valid_0 ? _GEN_96 : mask_0_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1121 = line_mask_clean_valid_0 ? _GEN_97 : mask_1_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1122 = line_mask_clean_valid_0 ? _GEN_98 : mask_2_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1123 = line_mask_clean_valid_0 ? _GEN_99 : mask_3_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1124 = line_mask_clean_valid_0 ? _GEN_100 : mask_4_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1125 = line_mask_clean_valid_0 ? _GEN_101 : mask_5_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1126 = line_mask_clean_valid_0 ? _GEN_102 : mask_6_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1127 = line_mask_clean_valid_0 ? _GEN_103 : mask_7_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1128 = line_mask_clean_valid_0 ? _GEN_104 : mask_8_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1129 = line_mask_clean_valid_0 ? _GEN_105 : mask_9_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1130 = line_mask_clean_valid_0 ? _GEN_106 : mask_10_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1131 = line_mask_clean_valid_0 ? _GEN_107 : mask_11_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1132 = line_mask_clean_valid_0 ? _GEN_108 : mask_12_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1133 = line_mask_clean_valid_0 ? _GEN_109 : mask_13_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1134 = line_mask_clean_valid_0 ? _GEN_110 : mask_14_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1135 = line_mask_clean_valid_0 ? _GEN_111 : mask_15_0_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1136 = line_mask_clean_valid_0 ? _GEN_112 : mask_0_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1137 = line_mask_clean_valid_0 ? _GEN_113 : mask_1_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1138 = line_mask_clean_valid_0 ? _GEN_114 : mask_2_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1139 = line_mask_clean_valid_0 ? _GEN_115 : mask_3_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1140 = line_mask_clean_valid_0 ? _GEN_116 : mask_4_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1141 = line_mask_clean_valid_0 ? _GEN_117 : mask_5_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1142 = line_mask_clean_valid_0 ? _GEN_118 : mask_6_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1143 = line_mask_clean_valid_0 ? _GEN_119 : mask_7_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1144 = line_mask_clean_valid_0 ? _GEN_120 : mask_8_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1145 = line_mask_clean_valid_0 ? _GEN_121 : mask_9_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1146 = line_mask_clean_valid_0 ? _GEN_122 : mask_10_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1147 = line_mask_clean_valid_0 ? _GEN_123 : mask_11_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1148 = line_mask_clean_valid_0 ? _GEN_124 : mask_12_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1149 = line_mask_clean_valid_0 ? _GEN_125 : mask_13_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1150 = line_mask_clean_valid_0 ? _GEN_126 : mask_14_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1151 = line_mask_clean_valid_0 ? _GEN_127 : mask_15_0_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1152 = line_mask_clean_valid_0 ? _GEN_128 : mask_0_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1153 = line_mask_clean_valid_0 ? _GEN_129 : mask_1_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1154 = line_mask_clean_valid_0 ? _GEN_130 : mask_2_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1155 = line_mask_clean_valid_0 ? _GEN_131 : mask_3_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1156 = line_mask_clean_valid_0 ? _GEN_132 : mask_4_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1157 = line_mask_clean_valid_0 ? _GEN_133 : mask_5_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1158 = line_mask_clean_valid_0 ? _GEN_134 : mask_6_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1159 = line_mask_clean_valid_0 ? _GEN_135 : mask_7_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1160 = line_mask_clean_valid_0 ? _GEN_136 : mask_8_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1161 = line_mask_clean_valid_0 ? _GEN_137 : mask_9_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1162 = line_mask_clean_valid_0 ? _GEN_138 : mask_10_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1163 = line_mask_clean_valid_0 ? _GEN_139 : mask_11_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1164 = line_mask_clean_valid_0 ? _GEN_140 : mask_12_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1165 = line_mask_clean_valid_0 ? _GEN_141 : mask_13_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1166 = line_mask_clean_valid_0 ? _GEN_142 : mask_14_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1167 = line_mask_clean_valid_0 ? _GEN_143 : mask_15_1_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1168 = line_mask_clean_valid_0 ? _GEN_144 : mask_0_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1169 = line_mask_clean_valid_0 ? _GEN_145 : mask_1_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1170 = line_mask_clean_valid_0 ? _GEN_146 : mask_2_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1171 = line_mask_clean_valid_0 ? _GEN_147 : mask_3_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1172 = line_mask_clean_valid_0 ? _GEN_148 : mask_4_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1173 = line_mask_clean_valid_0 ? _GEN_149 : mask_5_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1174 = line_mask_clean_valid_0 ? _GEN_150 : mask_6_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1175 = line_mask_clean_valid_0 ? _GEN_151 : mask_7_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1176 = line_mask_clean_valid_0 ? _GEN_152 : mask_8_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1177 = line_mask_clean_valid_0 ? _GEN_153 : mask_9_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1178 = line_mask_clean_valid_0 ? _GEN_154 : mask_10_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1179 = line_mask_clean_valid_0 ? _GEN_155 : mask_11_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1180 = line_mask_clean_valid_0 ? _GEN_156 : mask_12_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1181 = line_mask_clean_valid_0 ? _GEN_157 : mask_13_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1182 = line_mask_clean_valid_0 ? _GEN_158 : mask_14_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1183 = line_mask_clean_valid_0 ? _GEN_159 : mask_15_1_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1184 = line_mask_clean_valid_0 ? _GEN_160 : mask_0_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1185 = line_mask_clean_valid_0 ? _GEN_161 : mask_1_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1186 = line_mask_clean_valid_0 ? _GEN_162 : mask_2_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1187 = line_mask_clean_valid_0 ? _GEN_163 : mask_3_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1188 = line_mask_clean_valid_0 ? _GEN_164 : mask_4_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1189 = line_mask_clean_valid_0 ? _GEN_165 : mask_5_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1190 = line_mask_clean_valid_0 ? _GEN_166 : mask_6_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1191 = line_mask_clean_valid_0 ? _GEN_167 : mask_7_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1192 = line_mask_clean_valid_0 ? _GEN_168 : mask_8_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1193 = line_mask_clean_valid_0 ? _GEN_169 : mask_9_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1194 = line_mask_clean_valid_0 ? _GEN_170 : mask_10_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1195 = line_mask_clean_valid_0 ? _GEN_171 : mask_11_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1196 = line_mask_clean_valid_0 ? _GEN_172 : mask_12_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1197 = line_mask_clean_valid_0 ? _GEN_173 : mask_13_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1198 = line_mask_clean_valid_0 ? _GEN_174 : mask_14_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1199 = line_mask_clean_valid_0 ? _GEN_175 : mask_15_1_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1200 = line_mask_clean_valid_0 ? _GEN_176 : mask_0_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1201 = line_mask_clean_valid_0 ? _GEN_177 : mask_1_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1202 = line_mask_clean_valid_0 ? _GEN_178 : mask_2_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1203 = line_mask_clean_valid_0 ? _GEN_179 : mask_3_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1204 = line_mask_clean_valid_0 ? _GEN_180 : mask_4_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1205 = line_mask_clean_valid_0 ? _GEN_181 : mask_5_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1206 = line_mask_clean_valid_0 ? _GEN_182 : mask_6_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1207 = line_mask_clean_valid_0 ? _GEN_183 : mask_7_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1208 = line_mask_clean_valid_0 ? _GEN_184 : mask_8_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1209 = line_mask_clean_valid_0 ? _GEN_185 : mask_9_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1210 = line_mask_clean_valid_0 ? _GEN_186 : mask_10_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1211 = line_mask_clean_valid_0 ? _GEN_187 : mask_11_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1212 = line_mask_clean_valid_0 ? _GEN_188 : mask_12_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1213 = line_mask_clean_valid_0 ? _GEN_189 : mask_13_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1214 = line_mask_clean_valid_0 ? _GEN_190 : mask_14_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1215 = line_mask_clean_valid_0 ? _GEN_191 : mask_15_1_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1216 = line_mask_clean_valid_0 ? _GEN_192 : mask_0_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1217 = line_mask_clean_valid_0 ? _GEN_193 : mask_1_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1218 = line_mask_clean_valid_0 ? _GEN_194 : mask_2_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1219 = line_mask_clean_valid_0 ? _GEN_195 : mask_3_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1220 = line_mask_clean_valid_0 ? _GEN_196 : mask_4_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1221 = line_mask_clean_valid_0 ? _GEN_197 : mask_5_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1222 = line_mask_clean_valid_0 ? _GEN_198 : mask_6_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1223 = line_mask_clean_valid_0 ? _GEN_199 : mask_7_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1224 = line_mask_clean_valid_0 ? _GEN_200 : mask_8_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1225 = line_mask_clean_valid_0 ? _GEN_201 : mask_9_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1226 = line_mask_clean_valid_0 ? _GEN_202 : mask_10_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1227 = line_mask_clean_valid_0 ? _GEN_203 : mask_11_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1228 = line_mask_clean_valid_0 ? _GEN_204 : mask_12_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1229 = line_mask_clean_valid_0 ? _GEN_205 : mask_13_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1230 = line_mask_clean_valid_0 ? _GEN_206 : mask_14_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1231 = line_mask_clean_valid_0 ? _GEN_207 : mask_15_1_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1232 = line_mask_clean_valid_0 ? _GEN_208 : mask_0_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1233 = line_mask_clean_valid_0 ? _GEN_209 : mask_1_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1234 = line_mask_clean_valid_0 ? _GEN_210 : mask_2_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1235 = line_mask_clean_valid_0 ? _GEN_211 : mask_3_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1236 = line_mask_clean_valid_0 ? _GEN_212 : mask_4_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1237 = line_mask_clean_valid_0 ? _GEN_213 : mask_5_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1238 = line_mask_clean_valid_0 ? _GEN_214 : mask_6_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1239 = line_mask_clean_valid_0 ? _GEN_215 : mask_7_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1240 = line_mask_clean_valid_0 ? _GEN_216 : mask_8_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1241 = line_mask_clean_valid_0 ? _GEN_217 : mask_9_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1242 = line_mask_clean_valid_0 ? _GEN_218 : mask_10_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1243 = line_mask_clean_valid_0 ? _GEN_219 : mask_11_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1244 = line_mask_clean_valid_0 ? _GEN_220 : mask_12_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1245 = line_mask_clean_valid_0 ? _GEN_221 : mask_13_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1246 = line_mask_clean_valid_0 ? _GEN_222 : mask_14_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1247 = line_mask_clean_valid_0 ? _GEN_223 : mask_15_1_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1248 = line_mask_clean_valid_0 ? _GEN_224 : mask_0_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1249 = line_mask_clean_valid_0 ? _GEN_225 : mask_1_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1250 = line_mask_clean_valid_0 ? _GEN_226 : mask_2_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1251 = line_mask_clean_valid_0 ? _GEN_227 : mask_3_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1252 = line_mask_clean_valid_0 ? _GEN_228 : mask_4_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1253 = line_mask_clean_valid_0 ? _GEN_229 : mask_5_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1254 = line_mask_clean_valid_0 ? _GEN_230 : mask_6_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1255 = line_mask_clean_valid_0 ? _GEN_231 : mask_7_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1256 = line_mask_clean_valid_0 ? _GEN_232 : mask_8_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1257 = line_mask_clean_valid_0 ? _GEN_233 : mask_9_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1258 = line_mask_clean_valid_0 ? _GEN_234 : mask_10_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1259 = line_mask_clean_valid_0 ? _GEN_235 : mask_11_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1260 = line_mask_clean_valid_0 ? _GEN_236 : mask_12_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1261 = line_mask_clean_valid_0 ? _GEN_237 : mask_13_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1262 = line_mask_clean_valid_0 ? _GEN_238 : mask_14_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1263 = line_mask_clean_valid_0 ? _GEN_239 : mask_15_1_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1264 = line_mask_clean_valid_0 ? _GEN_240 : mask_0_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1265 = line_mask_clean_valid_0 ? _GEN_241 : mask_1_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1266 = line_mask_clean_valid_0 ? _GEN_242 : mask_2_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1267 = line_mask_clean_valid_0 ? _GEN_243 : mask_3_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1268 = line_mask_clean_valid_0 ? _GEN_244 : mask_4_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1269 = line_mask_clean_valid_0 ? _GEN_245 : mask_5_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1270 = line_mask_clean_valid_0 ? _GEN_246 : mask_6_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1271 = line_mask_clean_valid_0 ? _GEN_247 : mask_7_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1272 = line_mask_clean_valid_0 ? _GEN_248 : mask_8_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1273 = line_mask_clean_valid_0 ? _GEN_249 : mask_9_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1274 = line_mask_clean_valid_0 ? _GEN_250 : mask_10_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1275 = line_mask_clean_valid_0 ? _GEN_251 : mask_11_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1276 = line_mask_clean_valid_0 ? _GEN_252 : mask_12_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1277 = line_mask_clean_valid_0 ? _GEN_253 : mask_13_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1278 = line_mask_clean_valid_0 ? _GEN_254 : mask_14_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1279 = line_mask_clean_valid_0 ? _GEN_255 : mask_15_1_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1280 = line_mask_clean_valid_0 ? _GEN_256 : mask_0_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1281 = line_mask_clean_valid_0 ? _GEN_257 : mask_1_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1282 = line_mask_clean_valid_0 ? _GEN_258 : mask_2_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1283 = line_mask_clean_valid_0 ? _GEN_259 : mask_3_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1284 = line_mask_clean_valid_0 ? _GEN_260 : mask_4_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1285 = line_mask_clean_valid_0 ? _GEN_261 : mask_5_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1286 = line_mask_clean_valid_0 ? _GEN_262 : mask_6_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1287 = line_mask_clean_valid_0 ? _GEN_263 : mask_7_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1288 = line_mask_clean_valid_0 ? _GEN_264 : mask_8_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1289 = line_mask_clean_valid_0 ? _GEN_265 : mask_9_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1290 = line_mask_clean_valid_0 ? _GEN_266 : mask_10_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1291 = line_mask_clean_valid_0 ? _GEN_267 : mask_11_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1292 = line_mask_clean_valid_0 ? _GEN_268 : mask_12_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1293 = line_mask_clean_valid_0 ? _GEN_269 : mask_13_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1294 = line_mask_clean_valid_0 ? _GEN_270 : mask_14_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1295 = line_mask_clean_valid_0 ? _GEN_271 : mask_15_2_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1296 = line_mask_clean_valid_0 ? _GEN_272 : mask_0_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1297 = line_mask_clean_valid_0 ? _GEN_273 : mask_1_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1298 = line_mask_clean_valid_0 ? _GEN_274 : mask_2_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1299 = line_mask_clean_valid_0 ? _GEN_275 : mask_3_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1300 = line_mask_clean_valid_0 ? _GEN_276 : mask_4_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1301 = line_mask_clean_valid_0 ? _GEN_277 : mask_5_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1302 = line_mask_clean_valid_0 ? _GEN_278 : mask_6_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1303 = line_mask_clean_valid_0 ? _GEN_279 : mask_7_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1304 = line_mask_clean_valid_0 ? _GEN_280 : mask_8_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1305 = line_mask_clean_valid_0 ? _GEN_281 : mask_9_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1306 = line_mask_clean_valid_0 ? _GEN_282 : mask_10_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1307 = line_mask_clean_valid_0 ? _GEN_283 : mask_11_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1308 = line_mask_clean_valid_0 ? _GEN_284 : mask_12_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1309 = line_mask_clean_valid_0 ? _GEN_285 : mask_13_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1310 = line_mask_clean_valid_0 ? _GEN_286 : mask_14_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1311 = line_mask_clean_valid_0 ? _GEN_287 : mask_15_2_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1312 = line_mask_clean_valid_0 ? _GEN_288 : mask_0_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1313 = line_mask_clean_valid_0 ? _GEN_289 : mask_1_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1314 = line_mask_clean_valid_0 ? _GEN_290 : mask_2_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1315 = line_mask_clean_valid_0 ? _GEN_291 : mask_3_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1316 = line_mask_clean_valid_0 ? _GEN_292 : mask_4_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1317 = line_mask_clean_valid_0 ? _GEN_293 : mask_5_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1318 = line_mask_clean_valid_0 ? _GEN_294 : mask_6_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1319 = line_mask_clean_valid_0 ? _GEN_295 : mask_7_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1320 = line_mask_clean_valid_0 ? _GEN_296 : mask_8_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1321 = line_mask_clean_valid_0 ? _GEN_297 : mask_9_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1322 = line_mask_clean_valid_0 ? _GEN_298 : mask_10_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1323 = line_mask_clean_valid_0 ? _GEN_299 : mask_11_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1324 = line_mask_clean_valid_0 ? _GEN_300 : mask_12_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1325 = line_mask_clean_valid_0 ? _GEN_301 : mask_13_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1326 = line_mask_clean_valid_0 ? _GEN_302 : mask_14_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1327 = line_mask_clean_valid_0 ? _GEN_303 : mask_15_2_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1328 = line_mask_clean_valid_0 ? _GEN_304 : mask_0_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1329 = line_mask_clean_valid_0 ? _GEN_305 : mask_1_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1330 = line_mask_clean_valid_0 ? _GEN_306 : mask_2_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1331 = line_mask_clean_valid_0 ? _GEN_307 : mask_3_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1332 = line_mask_clean_valid_0 ? _GEN_308 : mask_4_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1333 = line_mask_clean_valid_0 ? _GEN_309 : mask_5_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1334 = line_mask_clean_valid_0 ? _GEN_310 : mask_6_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1335 = line_mask_clean_valid_0 ? _GEN_311 : mask_7_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1336 = line_mask_clean_valid_0 ? _GEN_312 : mask_8_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1337 = line_mask_clean_valid_0 ? _GEN_313 : mask_9_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1338 = line_mask_clean_valid_0 ? _GEN_314 : mask_10_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1339 = line_mask_clean_valid_0 ? _GEN_315 : mask_11_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1340 = line_mask_clean_valid_0 ? _GEN_316 : mask_12_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1341 = line_mask_clean_valid_0 ? _GEN_317 : mask_13_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1342 = line_mask_clean_valid_0 ? _GEN_318 : mask_14_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1343 = line_mask_clean_valid_0 ? _GEN_319 : mask_15_2_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1344 = line_mask_clean_valid_0 ? _GEN_320 : mask_0_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1345 = line_mask_clean_valid_0 ? _GEN_321 : mask_1_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1346 = line_mask_clean_valid_0 ? _GEN_322 : mask_2_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1347 = line_mask_clean_valid_0 ? _GEN_323 : mask_3_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1348 = line_mask_clean_valid_0 ? _GEN_324 : mask_4_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1349 = line_mask_clean_valid_0 ? _GEN_325 : mask_5_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1350 = line_mask_clean_valid_0 ? _GEN_326 : mask_6_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1351 = line_mask_clean_valid_0 ? _GEN_327 : mask_7_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1352 = line_mask_clean_valid_0 ? _GEN_328 : mask_8_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1353 = line_mask_clean_valid_0 ? _GEN_329 : mask_9_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1354 = line_mask_clean_valid_0 ? _GEN_330 : mask_10_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1355 = line_mask_clean_valid_0 ? _GEN_331 : mask_11_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1356 = line_mask_clean_valid_0 ? _GEN_332 : mask_12_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1357 = line_mask_clean_valid_0 ? _GEN_333 : mask_13_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1358 = line_mask_clean_valid_0 ? _GEN_334 : mask_14_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1359 = line_mask_clean_valid_0 ? _GEN_335 : mask_15_2_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1360 = line_mask_clean_valid_0 ? _GEN_336 : mask_0_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1361 = line_mask_clean_valid_0 ? _GEN_337 : mask_1_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1362 = line_mask_clean_valid_0 ? _GEN_338 : mask_2_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1363 = line_mask_clean_valid_0 ? _GEN_339 : mask_3_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1364 = line_mask_clean_valid_0 ? _GEN_340 : mask_4_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1365 = line_mask_clean_valid_0 ? _GEN_341 : mask_5_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1366 = line_mask_clean_valid_0 ? _GEN_342 : mask_6_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1367 = line_mask_clean_valid_0 ? _GEN_343 : mask_7_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1368 = line_mask_clean_valid_0 ? _GEN_344 : mask_8_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1369 = line_mask_clean_valid_0 ? _GEN_345 : mask_9_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1370 = line_mask_clean_valid_0 ? _GEN_346 : mask_10_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1371 = line_mask_clean_valid_0 ? _GEN_347 : mask_11_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1372 = line_mask_clean_valid_0 ? _GEN_348 : mask_12_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1373 = line_mask_clean_valid_0 ? _GEN_349 : mask_13_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1374 = line_mask_clean_valid_0 ? _GEN_350 : mask_14_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1375 = line_mask_clean_valid_0 ? _GEN_351 : mask_15_2_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1376 = line_mask_clean_valid_0 ? _GEN_352 : mask_0_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1377 = line_mask_clean_valid_0 ? _GEN_353 : mask_1_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1378 = line_mask_clean_valid_0 ? _GEN_354 : mask_2_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1379 = line_mask_clean_valid_0 ? _GEN_355 : mask_3_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1380 = line_mask_clean_valid_0 ? _GEN_356 : mask_4_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1381 = line_mask_clean_valid_0 ? _GEN_357 : mask_5_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1382 = line_mask_clean_valid_0 ? _GEN_358 : mask_6_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1383 = line_mask_clean_valid_0 ? _GEN_359 : mask_7_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1384 = line_mask_clean_valid_0 ? _GEN_360 : mask_8_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1385 = line_mask_clean_valid_0 ? _GEN_361 : mask_9_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1386 = line_mask_clean_valid_0 ? _GEN_362 : mask_10_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1387 = line_mask_clean_valid_0 ? _GEN_363 : mask_11_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1388 = line_mask_clean_valid_0 ? _GEN_364 : mask_12_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1389 = line_mask_clean_valid_0 ? _GEN_365 : mask_13_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1390 = line_mask_clean_valid_0 ? _GEN_366 : mask_14_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1391 = line_mask_clean_valid_0 ? _GEN_367 : mask_15_2_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1392 = line_mask_clean_valid_0 ? _GEN_368 : mask_0_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1393 = line_mask_clean_valid_0 ? _GEN_369 : mask_1_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1394 = line_mask_clean_valid_0 ? _GEN_370 : mask_2_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1395 = line_mask_clean_valid_0 ? _GEN_371 : mask_3_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1396 = line_mask_clean_valid_0 ? _GEN_372 : mask_4_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1397 = line_mask_clean_valid_0 ? _GEN_373 : mask_5_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1398 = line_mask_clean_valid_0 ? _GEN_374 : mask_6_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1399 = line_mask_clean_valid_0 ? _GEN_375 : mask_7_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1400 = line_mask_clean_valid_0 ? _GEN_376 : mask_8_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1401 = line_mask_clean_valid_0 ? _GEN_377 : mask_9_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1402 = line_mask_clean_valid_0 ? _GEN_378 : mask_10_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1403 = line_mask_clean_valid_0 ? _GEN_379 : mask_11_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1404 = line_mask_clean_valid_0 ? _GEN_380 : mask_12_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1405 = line_mask_clean_valid_0 ? _GEN_381 : mask_13_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1406 = line_mask_clean_valid_0 ? _GEN_382 : mask_14_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1407 = line_mask_clean_valid_0 ? _GEN_383 : mask_15_2_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1408 = line_mask_clean_valid_0 ? _GEN_384 : mask_0_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1409 = line_mask_clean_valid_0 ? _GEN_385 : mask_1_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1410 = line_mask_clean_valid_0 ? _GEN_386 : mask_2_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1411 = line_mask_clean_valid_0 ? _GEN_387 : mask_3_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1412 = line_mask_clean_valid_0 ? _GEN_388 : mask_4_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1413 = line_mask_clean_valid_0 ? _GEN_389 : mask_5_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1414 = line_mask_clean_valid_0 ? _GEN_390 : mask_6_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1415 = line_mask_clean_valid_0 ? _GEN_391 : mask_7_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1416 = line_mask_clean_valid_0 ? _GEN_392 : mask_8_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1417 = line_mask_clean_valid_0 ? _GEN_393 : mask_9_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1418 = line_mask_clean_valid_0 ? _GEN_394 : mask_10_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1419 = line_mask_clean_valid_0 ? _GEN_395 : mask_11_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1420 = line_mask_clean_valid_0 ? _GEN_396 : mask_12_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1421 = line_mask_clean_valid_0 ? _GEN_397 : mask_13_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1422 = line_mask_clean_valid_0 ? _GEN_398 : mask_14_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1423 = line_mask_clean_valid_0 ? _GEN_399 : mask_15_3_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1424 = line_mask_clean_valid_0 ? _GEN_400 : mask_0_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1425 = line_mask_clean_valid_0 ? _GEN_401 : mask_1_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1426 = line_mask_clean_valid_0 ? _GEN_402 : mask_2_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1427 = line_mask_clean_valid_0 ? _GEN_403 : mask_3_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1428 = line_mask_clean_valid_0 ? _GEN_404 : mask_4_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1429 = line_mask_clean_valid_0 ? _GEN_405 : mask_5_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1430 = line_mask_clean_valid_0 ? _GEN_406 : mask_6_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1431 = line_mask_clean_valid_0 ? _GEN_407 : mask_7_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1432 = line_mask_clean_valid_0 ? _GEN_408 : mask_8_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1433 = line_mask_clean_valid_0 ? _GEN_409 : mask_9_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1434 = line_mask_clean_valid_0 ? _GEN_410 : mask_10_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1435 = line_mask_clean_valid_0 ? _GEN_411 : mask_11_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1436 = line_mask_clean_valid_0 ? _GEN_412 : mask_12_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1437 = line_mask_clean_valid_0 ? _GEN_413 : mask_13_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1438 = line_mask_clean_valid_0 ? _GEN_414 : mask_14_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1439 = line_mask_clean_valid_0 ? _GEN_415 : mask_15_3_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1440 = line_mask_clean_valid_0 ? _GEN_416 : mask_0_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1441 = line_mask_clean_valid_0 ? _GEN_417 : mask_1_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1442 = line_mask_clean_valid_0 ? _GEN_418 : mask_2_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1443 = line_mask_clean_valid_0 ? _GEN_419 : mask_3_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1444 = line_mask_clean_valid_0 ? _GEN_420 : mask_4_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1445 = line_mask_clean_valid_0 ? _GEN_421 : mask_5_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1446 = line_mask_clean_valid_0 ? _GEN_422 : mask_6_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1447 = line_mask_clean_valid_0 ? _GEN_423 : mask_7_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1448 = line_mask_clean_valid_0 ? _GEN_424 : mask_8_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1449 = line_mask_clean_valid_0 ? _GEN_425 : mask_9_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1450 = line_mask_clean_valid_0 ? _GEN_426 : mask_10_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1451 = line_mask_clean_valid_0 ? _GEN_427 : mask_11_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1452 = line_mask_clean_valid_0 ? _GEN_428 : mask_12_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1453 = line_mask_clean_valid_0 ? _GEN_429 : mask_13_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1454 = line_mask_clean_valid_0 ? _GEN_430 : mask_14_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1455 = line_mask_clean_valid_0 ? _GEN_431 : mask_15_3_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1456 = line_mask_clean_valid_0 ? _GEN_432 : mask_0_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1457 = line_mask_clean_valid_0 ? _GEN_433 : mask_1_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1458 = line_mask_clean_valid_0 ? _GEN_434 : mask_2_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1459 = line_mask_clean_valid_0 ? _GEN_435 : mask_3_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1460 = line_mask_clean_valid_0 ? _GEN_436 : mask_4_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1461 = line_mask_clean_valid_0 ? _GEN_437 : mask_5_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1462 = line_mask_clean_valid_0 ? _GEN_438 : mask_6_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1463 = line_mask_clean_valid_0 ? _GEN_439 : mask_7_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1464 = line_mask_clean_valid_0 ? _GEN_440 : mask_8_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1465 = line_mask_clean_valid_0 ? _GEN_441 : mask_9_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1466 = line_mask_clean_valid_0 ? _GEN_442 : mask_10_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1467 = line_mask_clean_valid_0 ? _GEN_443 : mask_11_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1468 = line_mask_clean_valid_0 ? _GEN_444 : mask_12_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1469 = line_mask_clean_valid_0 ? _GEN_445 : mask_13_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1470 = line_mask_clean_valid_0 ? _GEN_446 : mask_14_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1471 = line_mask_clean_valid_0 ? _GEN_447 : mask_15_3_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1472 = line_mask_clean_valid_0 ? _GEN_448 : mask_0_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1473 = line_mask_clean_valid_0 ? _GEN_449 : mask_1_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1474 = line_mask_clean_valid_0 ? _GEN_450 : mask_2_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1475 = line_mask_clean_valid_0 ? _GEN_451 : mask_3_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1476 = line_mask_clean_valid_0 ? _GEN_452 : mask_4_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1477 = line_mask_clean_valid_0 ? _GEN_453 : mask_5_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1478 = line_mask_clean_valid_0 ? _GEN_454 : mask_6_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1479 = line_mask_clean_valid_0 ? _GEN_455 : mask_7_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1480 = line_mask_clean_valid_0 ? _GEN_456 : mask_8_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1481 = line_mask_clean_valid_0 ? _GEN_457 : mask_9_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1482 = line_mask_clean_valid_0 ? _GEN_458 : mask_10_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1483 = line_mask_clean_valid_0 ? _GEN_459 : mask_11_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1484 = line_mask_clean_valid_0 ? _GEN_460 : mask_12_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1485 = line_mask_clean_valid_0 ? _GEN_461 : mask_13_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1486 = line_mask_clean_valid_0 ? _GEN_462 : mask_14_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1487 = line_mask_clean_valid_0 ? _GEN_463 : mask_15_3_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1488 = line_mask_clean_valid_0 ? _GEN_464 : mask_0_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1489 = line_mask_clean_valid_0 ? _GEN_465 : mask_1_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1490 = line_mask_clean_valid_0 ? _GEN_466 : mask_2_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1491 = line_mask_clean_valid_0 ? _GEN_467 : mask_3_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1492 = line_mask_clean_valid_0 ? _GEN_468 : mask_4_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1493 = line_mask_clean_valid_0 ? _GEN_469 : mask_5_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1494 = line_mask_clean_valid_0 ? _GEN_470 : mask_6_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1495 = line_mask_clean_valid_0 ? _GEN_471 : mask_7_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1496 = line_mask_clean_valid_0 ? _GEN_472 : mask_8_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1497 = line_mask_clean_valid_0 ? _GEN_473 : mask_9_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1498 = line_mask_clean_valid_0 ? _GEN_474 : mask_10_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1499 = line_mask_clean_valid_0 ? _GEN_475 : mask_11_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1500 = line_mask_clean_valid_0 ? _GEN_476 : mask_12_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1501 = line_mask_clean_valid_0 ? _GEN_477 : mask_13_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1502 = line_mask_clean_valid_0 ? _GEN_478 : mask_14_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1503 = line_mask_clean_valid_0 ? _GEN_479 : mask_15_3_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1504 = line_mask_clean_valid_0 ? _GEN_480 : mask_0_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1505 = line_mask_clean_valid_0 ? _GEN_481 : mask_1_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1506 = line_mask_clean_valid_0 ? _GEN_482 : mask_2_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1507 = line_mask_clean_valid_0 ? _GEN_483 : mask_3_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1508 = line_mask_clean_valid_0 ? _GEN_484 : mask_4_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1509 = line_mask_clean_valid_0 ? _GEN_485 : mask_5_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1510 = line_mask_clean_valid_0 ? _GEN_486 : mask_6_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1511 = line_mask_clean_valid_0 ? _GEN_487 : mask_7_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1512 = line_mask_clean_valid_0 ? _GEN_488 : mask_8_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1513 = line_mask_clean_valid_0 ? _GEN_489 : mask_9_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1514 = line_mask_clean_valid_0 ? _GEN_490 : mask_10_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1515 = line_mask_clean_valid_0 ? _GEN_491 : mask_11_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1516 = line_mask_clean_valid_0 ? _GEN_492 : mask_12_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1517 = line_mask_clean_valid_0 ? _GEN_493 : mask_13_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1518 = line_mask_clean_valid_0 ? _GEN_494 : mask_14_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1519 = line_mask_clean_valid_0 ? _GEN_495 : mask_15_3_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1520 = line_mask_clean_valid_0 ? _GEN_496 : mask_0_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1521 = line_mask_clean_valid_0 ? _GEN_497 : mask_1_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1522 = line_mask_clean_valid_0 ? _GEN_498 : mask_2_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1523 = line_mask_clean_valid_0 ? _GEN_499 : mask_3_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1524 = line_mask_clean_valid_0 ? _GEN_500 : mask_4_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1525 = line_mask_clean_valid_0 ? _GEN_501 : mask_5_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1526 = line_mask_clean_valid_0 ? _GEN_502 : mask_6_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1527 = line_mask_clean_valid_0 ? _GEN_503 : mask_7_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1528 = line_mask_clean_valid_0 ? _GEN_504 : mask_8_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1529 = line_mask_clean_valid_0 ? _GEN_505 : mask_9_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1530 = line_mask_clean_valid_0 ? _GEN_506 : mask_10_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1531 = line_mask_clean_valid_0 ? _GEN_507 : mask_11_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1532 = line_mask_clean_valid_0 ? _GEN_508 : mask_12_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1533 = line_mask_clean_valid_0 ? _GEN_509 : mask_13_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1534 = line_mask_clean_valid_0 ? _GEN_510 : mask_14_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1535 = line_mask_clean_valid_0 ? _GEN_511 : mask_15_3_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1536 = line_mask_clean_valid_0 ? _GEN_512 : mask_0_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1537 = line_mask_clean_valid_0 ? _GEN_513 : mask_1_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1538 = line_mask_clean_valid_0 ? _GEN_514 : mask_2_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1539 = line_mask_clean_valid_0 ? _GEN_515 : mask_3_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1540 = line_mask_clean_valid_0 ? _GEN_516 : mask_4_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1541 = line_mask_clean_valid_0 ? _GEN_517 : mask_5_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1542 = line_mask_clean_valid_0 ? _GEN_518 : mask_6_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1543 = line_mask_clean_valid_0 ? _GEN_519 : mask_7_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1544 = line_mask_clean_valid_0 ? _GEN_520 : mask_8_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1545 = line_mask_clean_valid_0 ? _GEN_521 : mask_9_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1546 = line_mask_clean_valid_0 ? _GEN_522 : mask_10_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1547 = line_mask_clean_valid_0 ? _GEN_523 : mask_11_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1548 = line_mask_clean_valid_0 ? _GEN_524 : mask_12_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1549 = line_mask_clean_valid_0 ? _GEN_525 : mask_13_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1550 = line_mask_clean_valid_0 ? _GEN_526 : mask_14_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1551 = line_mask_clean_valid_0 ? _GEN_527 : mask_15_4_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1552 = line_mask_clean_valid_0 ? _GEN_528 : mask_0_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1553 = line_mask_clean_valid_0 ? _GEN_529 : mask_1_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1554 = line_mask_clean_valid_0 ? _GEN_530 : mask_2_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1555 = line_mask_clean_valid_0 ? _GEN_531 : mask_3_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1556 = line_mask_clean_valid_0 ? _GEN_532 : mask_4_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1557 = line_mask_clean_valid_0 ? _GEN_533 : mask_5_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1558 = line_mask_clean_valid_0 ? _GEN_534 : mask_6_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1559 = line_mask_clean_valid_0 ? _GEN_535 : mask_7_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1560 = line_mask_clean_valid_0 ? _GEN_536 : mask_8_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1561 = line_mask_clean_valid_0 ? _GEN_537 : mask_9_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1562 = line_mask_clean_valid_0 ? _GEN_538 : mask_10_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1563 = line_mask_clean_valid_0 ? _GEN_539 : mask_11_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1564 = line_mask_clean_valid_0 ? _GEN_540 : mask_12_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1565 = line_mask_clean_valid_0 ? _GEN_541 : mask_13_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1566 = line_mask_clean_valid_0 ? _GEN_542 : mask_14_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1567 = line_mask_clean_valid_0 ? _GEN_543 : mask_15_4_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1568 = line_mask_clean_valid_0 ? _GEN_544 : mask_0_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1569 = line_mask_clean_valid_0 ? _GEN_545 : mask_1_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1570 = line_mask_clean_valid_0 ? _GEN_546 : mask_2_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1571 = line_mask_clean_valid_0 ? _GEN_547 : mask_3_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1572 = line_mask_clean_valid_0 ? _GEN_548 : mask_4_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1573 = line_mask_clean_valid_0 ? _GEN_549 : mask_5_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1574 = line_mask_clean_valid_0 ? _GEN_550 : mask_6_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1575 = line_mask_clean_valid_0 ? _GEN_551 : mask_7_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1576 = line_mask_clean_valid_0 ? _GEN_552 : mask_8_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1577 = line_mask_clean_valid_0 ? _GEN_553 : mask_9_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1578 = line_mask_clean_valid_0 ? _GEN_554 : mask_10_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1579 = line_mask_clean_valid_0 ? _GEN_555 : mask_11_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1580 = line_mask_clean_valid_0 ? _GEN_556 : mask_12_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1581 = line_mask_clean_valid_0 ? _GEN_557 : mask_13_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1582 = line_mask_clean_valid_0 ? _GEN_558 : mask_14_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1583 = line_mask_clean_valid_0 ? _GEN_559 : mask_15_4_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1584 = line_mask_clean_valid_0 ? _GEN_560 : mask_0_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1585 = line_mask_clean_valid_0 ? _GEN_561 : mask_1_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1586 = line_mask_clean_valid_0 ? _GEN_562 : mask_2_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1587 = line_mask_clean_valid_0 ? _GEN_563 : mask_3_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1588 = line_mask_clean_valid_0 ? _GEN_564 : mask_4_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1589 = line_mask_clean_valid_0 ? _GEN_565 : mask_5_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1590 = line_mask_clean_valid_0 ? _GEN_566 : mask_6_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1591 = line_mask_clean_valid_0 ? _GEN_567 : mask_7_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1592 = line_mask_clean_valid_0 ? _GEN_568 : mask_8_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1593 = line_mask_clean_valid_0 ? _GEN_569 : mask_9_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1594 = line_mask_clean_valid_0 ? _GEN_570 : mask_10_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1595 = line_mask_clean_valid_0 ? _GEN_571 : mask_11_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1596 = line_mask_clean_valid_0 ? _GEN_572 : mask_12_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1597 = line_mask_clean_valid_0 ? _GEN_573 : mask_13_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1598 = line_mask_clean_valid_0 ? _GEN_574 : mask_14_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1599 = line_mask_clean_valid_0 ? _GEN_575 : mask_15_4_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1600 = line_mask_clean_valid_0 ? _GEN_576 : mask_0_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1601 = line_mask_clean_valid_0 ? _GEN_577 : mask_1_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1602 = line_mask_clean_valid_0 ? _GEN_578 : mask_2_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1603 = line_mask_clean_valid_0 ? _GEN_579 : mask_3_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1604 = line_mask_clean_valid_0 ? _GEN_580 : mask_4_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1605 = line_mask_clean_valid_0 ? _GEN_581 : mask_5_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1606 = line_mask_clean_valid_0 ? _GEN_582 : mask_6_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1607 = line_mask_clean_valid_0 ? _GEN_583 : mask_7_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1608 = line_mask_clean_valid_0 ? _GEN_584 : mask_8_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1609 = line_mask_clean_valid_0 ? _GEN_585 : mask_9_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1610 = line_mask_clean_valid_0 ? _GEN_586 : mask_10_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1611 = line_mask_clean_valid_0 ? _GEN_587 : mask_11_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1612 = line_mask_clean_valid_0 ? _GEN_588 : mask_12_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1613 = line_mask_clean_valid_0 ? _GEN_589 : mask_13_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1614 = line_mask_clean_valid_0 ? _GEN_590 : mask_14_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1615 = line_mask_clean_valid_0 ? _GEN_591 : mask_15_4_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1616 = line_mask_clean_valid_0 ? _GEN_592 : mask_0_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1617 = line_mask_clean_valid_0 ? _GEN_593 : mask_1_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1618 = line_mask_clean_valid_0 ? _GEN_594 : mask_2_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1619 = line_mask_clean_valid_0 ? _GEN_595 : mask_3_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1620 = line_mask_clean_valid_0 ? _GEN_596 : mask_4_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1621 = line_mask_clean_valid_0 ? _GEN_597 : mask_5_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1622 = line_mask_clean_valid_0 ? _GEN_598 : mask_6_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1623 = line_mask_clean_valid_0 ? _GEN_599 : mask_7_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1624 = line_mask_clean_valid_0 ? _GEN_600 : mask_8_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1625 = line_mask_clean_valid_0 ? _GEN_601 : mask_9_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1626 = line_mask_clean_valid_0 ? _GEN_602 : mask_10_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1627 = line_mask_clean_valid_0 ? _GEN_603 : mask_11_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1628 = line_mask_clean_valid_0 ? _GEN_604 : mask_12_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1629 = line_mask_clean_valid_0 ? _GEN_605 : mask_13_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1630 = line_mask_clean_valid_0 ? _GEN_606 : mask_14_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1631 = line_mask_clean_valid_0 ? _GEN_607 : mask_15_4_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1632 = line_mask_clean_valid_0 ? _GEN_608 : mask_0_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1633 = line_mask_clean_valid_0 ? _GEN_609 : mask_1_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1634 = line_mask_clean_valid_0 ? _GEN_610 : mask_2_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1635 = line_mask_clean_valid_0 ? _GEN_611 : mask_3_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1636 = line_mask_clean_valid_0 ? _GEN_612 : mask_4_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1637 = line_mask_clean_valid_0 ? _GEN_613 : mask_5_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1638 = line_mask_clean_valid_0 ? _GEN_614 : mask_6_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1639 = line_mask_clean_valid_0 ? _GEN_615 : mask_7_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1640 = line_mask_clean_valid_0 ? _GEN_616 : mask_8_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1641 = line_mask_clean_valid_0 ? _GEN_617 : mask_9_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1642 = line_mask_clean_valid_0 ? _GEN_618 : mask_10_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1643 = line_mask_clean_valid_0 ? _GEN_619 : mask_11_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1644 = line_mask_clean_valid_0 ? _GEN_620 : mask_12_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1645 = line_mask_clean_valid_0 ? _GEN_621 : mask_13_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1646 = line_mask_clean_valid_0 ? _GEN_622 : mask_14_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1647 = line_mask_clean_valid_0 ? _GEN_623 : mask_15_4_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1648 = line_mask_clean_valid_0 ? _GEN_624 : mask_0_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1649 = line_mask_clean_valid_0 ? _GEN_625 : mask_1_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1650 = line_mask_clean_valid_0 ? _GEN_626 : mask_2_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1651 = line_mask_clean_valid_0 ? _GEN_627 : mask_3_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1652 = line_mask_clean_valid_0 ? _GEN_628 : mask_4_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1653 = line_mask_clean_valid_0 ? _GEN_629 : mask_5_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1654 = line_mask_clean_valid_0 ? _GEN_630 : mask_6_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1655 = line_mask_clean_valid_0 ? _GEN_631 : mask_7_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1656 = line_mask_clean_valid_0 ? _GEN_632 : mask_8_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1657 = line_mask_clean_valid_0 ? _GEN_633 : mask_9_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1658 = line_mask_clean_valid_0 ? _GEN_634 : mask_10_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1659 = line_mask_clean_valid_0 ? _GEN_635 : mask_11_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1660 = line_mask_clean_valid_0 ? _GEN_636 : mask_12_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1661 = line_mask_clean_valid_0 ? _GEN_637 : mask_13_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1662 = line_mask_clean_valid_0 ? _GEN_638 : mask_14_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1663 = line_mask_clean_valid_0 ? _GEN_639 : mask_15_4_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1664 = line_mask_clean_valid_0 ? _GEN_640 : mask_0_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1665 = line_mask_clean_valid_0 ? _GEN_641 : mask_1_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1666 = line_mask_clean_valid_0 ? _GEN_642 : mask_2_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1667 = line_mask_clean_valid_0 ? _GEN_643 : mask_3_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1668 = line_mask_clean_valid_0 ? _GEN_644 : mask_4_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1669 = line_mask_clean_valid_0 ? _GEN_645 : mask_5_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1670 = line_mask_clean_valid_0 ? _GEN_646 : mask_6_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1671 = line_mask_clean_valid_0 ? _GEN_647 : mask_7_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1672 = line_mask_clean_valid_0 ? _GEN_648 : mask_8_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1673 = line_mask_clean_valid_0 ? _GEN_649 : mask_9_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1674 = line_mask_clean_valid_0 ? _GEN_650 : mask_10_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1675 = line_mask_clean_valid_0 ? _GEN_651 : mask_11_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1676 = line_mask_clean_valid_0 ? _GEN_652 : mask_12_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1677 = line_mask_clean_valid_0 ? _GEN_653 : mask_13_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1678 = line_mask_clean_valid_0 ? _GEN_654 : mask_14_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1679 = line_mask_clean_valid_0 ? _GEN_655 : mask_15_5_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1680 = line_mask_clean_valid_0 ? _GEN_656 : mask_0_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1681 = line_mask_clean_valid_0 ? _GEN_657 : mask_1_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1682 = line_mask_clean_valid_0 ? _GEN_658 : mask_2_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1683 = line_mask_clean_valid_0 ? _GEN_659 : mask_3_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1684 = line_mask_clean_valid_0 ? _GEN_660 : mask_4_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1685 = line_mask_clean_valid_0 ? _GEN_661 : mask_5_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1686 = line_mask_clean_valid_0 ? _GEN_662 : mask_6_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1687 = line_mask_clean_valid_0 ? _GEN_663 : mask_7_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1688 = line_mask_clean_valid_0 ? _GEN_664 : mask_8_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1689 = line_mask_clean_valid_0 ? _GEN_665 : mask_9_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1690 = line_mask_clean_valid_0 ? _GEN_666 : mask_10_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1691 = line_mask_clean_valid_0 ? _GEN_667 : mask_11_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1692 = line_mask_clean_valid_0 ? _GEN_668 : mask_12_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1693 = line_mask_clean_valid_0 ? _GEN_669 : mask_13_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1694 = line_mask_clean_valid_0 ? _GEN_670 : mask_14_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1695 = line_mask_clean_valid_0 ? _GEN_671 : mask_15_5_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1696 = line_mask_clean_valid_0 ? _GEN_672 : mask_0_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1697 = line_mask_clean_valid_0 ? _GEN_673 : mask_1_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1698 = line_mask_clean_valid_0 ? _GEN_674 : mask_2_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1699 = line_mask_clean_valid_0 ? _GEN_675 : mask_3_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1700 = line_mask_clean_valid_0 ? _GEN_676 : mask_4_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1701 = line_mask_clean_valid_0 ? _GEN_677 : mask_5_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1702 = line_mask_clean_valid_0 ? _GEN_678 : mask_6_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1703 = line_mask_clean_valid_0 ? _GEN_679 : mask_7_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1704 = line_mask_clean_valid_0 ? _GEN_680 : mask_8_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1705 = line_mask_clean_valid_0 ? _GEN_681 : mask_9_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1706 = line_mask_clean_valid_0 ? _GEN_682 : mask_10_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1707 = line_mask_clean_valid_0 ? _GEN_683 : mask_11_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1708 = line_mask_clean_valid_0 ? _GEN_684 : mask_12_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1709 = line_mask_clean_valid_0 ? _GEN_685 : mask_13_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1710 = line_mask_clean_valid_0 ? _GEN_686 : mask_14_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1711 = line_mask_clean_valid_0 ? _GEN_687 : mask_15_5_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1712 = line_mask_clean_valid_0 ? _GEN_688 : mask_0_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1713 = line_mask_clean_valid_0 ? _GEN_689 : mask_1_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1714 = line_mask_clean_valid_0 ? _GEN_690 : mask_2_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1715 = line_mask_clean_valid_0 ? _GEN_691 : mask_3_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1716 = line_mask_clean_valid_0 ? _GEN_692 : mask_4_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1717 = line_mask_clean_valid_0 ? _GEN_693 : mask_5_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1718 = line_mask_clean_valid_0 ? _GEN_694 : mask_6_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1719 = line_mask_clean_valid_0 ? _GEN_695 : mask_7_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1720 = line_mask_clean_valid_0 ? _GEN_696 : mask_8_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1721 = line_mask_clean_valid_0 ? _GEN_697 : mask_9_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1722 = line_mask_clean_valid_0 ? _GEN_698 : mask_10_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1723 = line_mask_clean_valid_0 ? _GEN_699 : mask_11_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1724 = line_mask_clean_valid_0 ? _GEN_700 : mask_12_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1725 = line_mask_clean_valid_0 ? _GEN_701 : mask_13_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1726 = line_mask_clean_valid_0 ? _GEN_702 : mask_14_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1727 = line_mask_clean_valid_0 ? _GEN_703 : mask_15_5_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1728 = line_mask_clean_valid_0 ? _GEN_704 : mask_0_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1729 = line_mask_clean_valid_0 ? _GEN_705 : mask_1_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1730 = line_mask_clean_valid_0 ? _GEN_706 : mask_2_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1731 = line_mask_clean_valid_0 ? _GEN_707 : mask_3_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1732 = line_mask_clean_valid_0 ? _GEN_708 : mask_4_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1733 = line_mask_clean_valid_0 ? _GEN_709 : mask_5_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1734 = line_mask_clean_valid_0 ? _GEN_710 : mask_6_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1735 = line_mask_clean_valid_0 ? _GEN_711 : mask_7_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1736 = line_mask_clean_valid_0 ? _GEN_712 : mask_8_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1737 = line_mask_clean_valid_0 ? _GEN_713 : mask_9_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1738 = line_mask_clean_valid_0 ? _GEN_714 : mask_10_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1739 = line_mask_clean_valid_0 ? _GEN_715 : mask_11_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1740 = line_mask_clean_valid_0 ? _GEN_716 : mask_12_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1741 = line_mask_clean_valid_0 ? _GEN_717 : mask_13_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1742 = line_mask_clean_valid_0 ? _GEN_718 : mask_14_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1743 = line_mask_clean_valid_0 ? _GEN_719 : mask_15_5_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1744 = line_mask_clean_valid_0 ? _GEN_720 : mask_0_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1745 = line_mask_clean_valid_0 ? _GEN_721 : mask_1_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1746 = line_mask_clean_valid_0 ? _GEN_722 : mask_2_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1747 = line_mask_clean_valid_0 ? _GEN_723 : mask_3_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1748 = line_mask_clean_valid_0 ? _GEN_724 : mask_4_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1749 = line_mask_clean_valid_0 ? _GEN_725 : mask_5_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1750 = line_mask_clean_valid_0 ? _GEN_726 : mask_6_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1751 = line_mask_clean_valid_0 ? _GEN_727 : mask_7_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1752 = line_mask_clean_valid_0 ? _GEN_728 : mask_8_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1753 = line_mask_clean_valid_0 ? _GEN_729 : mask_9_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1754 = line_mask_clean_valid_0 ? _GEN_730 : mask_10_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1755 = line_mask_clean_valid_0 ? _GEN_731 : mask_11_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1756 = line_mask_clean_valid_0 ? _GEN_732 : mask_12_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1757 = line_mask_clean_valid_0 ? _GEN_733 : mask_13_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1758 = line_mask_clean_valid_0 ? _GEN_734 : mask_14_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1759 = line_mask_clean_valid_0 ? _GEN_735 : mask_15_5_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1760 = line_mask_clean_valid_0 ? _GEN_736 : mask_0_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1761 = line_mask_clean_valid_0 ? _GEN_737 : mask_1_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1762 = line_mask_clean_valid_0 ? _GEN_738 : mask_2_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1763 = line_mask_clean_valid_0 ? _GEN_739 : mask_3_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1764 = line_mask_clean_valid_0 ? _GEN_740 : mask_4_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1765 = line_mask_clean_valid_0 ? _GEN_741 : mask_5_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1766 = line_mask_clean_valid_0 ? _GEN_742 : mask_6_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1767 = line_mask_clean_valid_0 ? _GEN_743 : mask_7_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1768 = line_mask_clean_valid_0 ? _GEN_744 : mask_8_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1769 = line_mask_clean_valid_0 ? _GEN_745 : mask_9_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1770 = line_mask_clean_valid_0 ? _GEN_746 : mask_10_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1771 = line_mask_clean_valid_0 ? _GEN_747 : mask_11_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1772 = line_mask_clean_valid_0 ? _GEN_748 : mask_12_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1773 = line_mask_clean_valid_0 ? _GEN_749 : mask_13_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1774 = line_mask_clean_valid_0 ? _GEN_750 : mask_14_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1775 = line_mask_clean_valid_0 ? _GEN_751 : mask_15_5_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1776 = line_mask_clean_valid_0 ? _GEN_752 : mask_0_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1777 = line_mask_clean_valid_0 ? _GEN_753 : mask_1_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1778 = line_mask_clean_valid_0 ? _GEN_754 : mask_2_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1779 = line_mask_clean_valid_0 ? _GEN_755 : mask_3_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1780 = line_mask_clean_valid_0 ? _GEN_756 : mask_4_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1781 = line_mask_clean_valid_0 ? _GEN_757 : mask_5_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1782 = line_mask_clean_valid_0 ? _GEN_758 : mask_6_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1783 = line_mask_clean_valid_0 ? _GEN_759 : mask_7_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1784 = line_mask_clean_valid_0 ? _GEN_760 : mask_8_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1785 = line_mask_clean_valid_0 ? _GEN_761 : mask_9_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1786 = line_mask_clean_valid_0 ? _GEN_762 : mask_10_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1787 = line_mask_clean_valid_0 ? _GEN_763 : mask_11_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1788 = line_mask_clean_valid_0 ? _GEN_764 : mask_12_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1789 = line_mask_clean_valid_0 ? _GEN_765 : mask_13_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1790 = line_mask_clean_valid_0 ? _GEN_766 : mask_14_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1791 = line_mask_clean_valid_0 ? _GEN_767 : mask_15_5_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1792 = line_mask_clean_valid_0 ? _GEN_768 : mask_0_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1793 = line_mask_clean_valid_0 ? _GEN_769 : mask_1_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1794 = line_mask_clean_valid_0 ? _GEN_770 : mask_2_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1795 = line_mask_clean_valid_0 ? _GEN_771 : mask_3_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1796 = line_mask_clean_valid_0 ? _GEN_772 : mask_4_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1797 = line_mask_clean_valid_0 ? _GEN_773 : mask_5_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1798 = line_mask_clean_valid_0 ? _GEN_774 : mask_6_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1799 = line_mask_clean_valid_0 ? _GEN_775 : mask_7_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1800 = line_mask_clean_valid_0 ? _GEN_776 : mask_8_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1801 = line_mask_clean_valid_0 ? _GEN_777 : mask_9_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1802 = line_mask_clean_valid_0 ? _GEN_778 : mask_10_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1803 = line_mask_clean_valid_0 ? _GEN_779 : mask_11_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1804 = line_mask_clean_valid_0 ? _GEN_780 : mask_12_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1805 = line_mask_clean_valid_0 ? _GEN_781 : mask_13_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1806 = line_mask_clean_valid_0 ? _GEN_782 : mask_14_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1807 = line_mask_clean_valid_0 ? _GEN_783 : mask_15_6_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1808 = line_mask_clean_valid_0 ? _GEN_784 : mask_0_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1809 = line_mask_clean_valid_0 ? _GEN_785 : mask_1_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1810 = line_mask_clean_valid_0 ? _GEN_786 : mask_2_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1811 = line_mask_clean_valid_0 ? _GEN_787 : mask_3_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1812 = line_mask_clean_valid_0 ? _GEN_788 : mask_4_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1813 = line_mask_clean_valid_0 ? _GEN_789 : mask_5_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1814 = line_mask_clean_valid_0 ? _GEN_790 : mask_6_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1815 = line_mask_clean_valid_0 ? _GEN_791 : mask_7_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1816 = line_mask_clean_valid_0 ? _GEN_792 : mask_8_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1817 = line_mask_clean_valid_0 ? _GEN_793 : mask_9_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1818 = line_mask_clean_valid_0 ? _GEN_794 : mask_10_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1819 = line_mask_clean_valid_0 ? _GEN_795 : mask_11_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1820 = line_mask_clean_valid_0 ? _GEN_796 : mask_12_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1821 = line_mask_clean_valid_0 ? _GEN_797 : mask_13_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1822 = line_mask_clean_valid_0 ? _GEN_798 : mask_14_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1823 = line_mask_clean_valid_0 ? _GEN_799 : mask_15_6_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1824 = line_mask_clean_valid_0 ? _GEN_800 : mask_0_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1825 = line_mask_clean_valid_0 ? _GEN_801 : mask_1_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1826 = line_mask_clean_valid_0 ? _GEN_802 : mask_2_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1827 = line_mask_clean_valid_0 ? _GEN_803 : mask_3_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1828 = line_mask_clean_valid_0 ? _GEN_804 : mask_4_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1829 = line_mask_clean_valid_0 ? _GEN_805 : mask_5_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1830 = line_mask_clean_valid_0 ? _GEN_806 : mask_6_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1831 = line_mask_clean_valid_0 ? _GEN_807 : mask_7_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1832 = line_mask_clean_valid_0 ? _GEN_808 : mask_8_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1833 = line_mask_clean_valid_0 ? _GEN_809 : mask_9_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1834 = line_mask_clean_valid_0 ? _GEN_810 : mask_10_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1835 = line_mask_clean_valid_0 ? _GEN_811 : mask_11_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1836 = line_mask_clean_valid_0 ? _GEN_812 : mask_12_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1837 = line_mask_clean_valid_0 ? _GEN_813 : mask_13_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1838 = line_mask_clean_valid_0 ? _GEN_814 : mask_14_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1839 = line_mask_clean_valid_0 ? _GEN_815 : mask_15_6_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1840 = line_mask_clean_valid_0 ? _GEN_816 : mask_0_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1841 = line_mask_clean_valid_0 ? _GEN_817 : mask_1_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1842 = line_mask_clean_valid_0 ? _GEN_818 : mask_2_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1843 = line_mask_clean_valid_0 ? _GEN_819 : mask_3_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1844 = line_mask_clean_valid_0 ? _GEN_820 : mask_4_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1845 = line_mask_clean_valid_0 ? _GEN_821 : mask_5_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1846 = line_mask_clean_valid_0 ? _GEN_822 : mask_6_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1847 = line_mask_clean_valid_0 ? _GEN_823 : mask_7_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1848 = line_mask_clean_valid_0 ? _GEN_824 : mask_8_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1849 = line_mask_clean_valid_0 ? _GEN_825 : mask_9_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1850 = line_mask_clean_valid_0 ? _GEN_826 : mask_10_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1851 = line_mask_clean_valid_0 ? _GEN_827 : mask_11_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1852 = line_mask_clean_valid_0 ? _GEN_828 : mask_12_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1853 = line_mask_clean_valid_0 ? _GEN_829 : mask_13_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1854 = line_mask_clean_valid_0 ? _GEN_830 : mask_14_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1855 = line_mask_clean_valid_0 ? _GEN_831 : mask_15_6_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1856 = line_mask_clean_valid_0 ? _GEN_832 : mask_0_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1857 = line_mask_clean_valid_0 ? _GEN_833 : mask_1_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1858 = line_mask_clean_valid_0 ? _GEN_834 : mask_2_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1859 = line_mask_clean_valid_0 ? _GEN_835 : mask_3_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1860 = line_mask_clean_valid_0 ? _GEN_836 : mask_4_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1861 = line_mask_clean_valid_0 ? _GEN_837 : mask_5_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1862 = line_mask_clean_valid_0 ? _GEN_838 : mask_6_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1863 = line_mask_clean_valid_0 ? _GEN_839 : mask_7_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1864 = line_mask_clean_valid_0 ? _GEN_840 : mask_8_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1865 = line_mask_clean_valid_0 ? _GEN_841 : mask_9_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1866 = line_mask_clean_valid_0 ? _GEN_842 : mask_10_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1867 = line_mask_clean_valid_0 ? _GEN_843 : mask_11_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1868 = line_mask_clean_valid_0 ? _GEN_844 : mask_12_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1869 = line_mask_clean_valid_0 ? _GEN_845 : mask_13_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1870 = line_mask_clean_valid_0 ? _GEN_846 : mask_14_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1871 = line_mask_clean_valid_0 ? _GEN_847 : mask_15_6_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1872 = line_mask_clean_valid_0 ? _GEN_848 : mask_0_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1873 = line_mask_clean_valid_0 ? _GEN_849 : mask_1_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1874 = line_mask_clean_valid_0 ? _GEN_850 : mask_2_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1875 = line_mask_clean_valid_0 ? _GEN_851 : mask_3_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1876 = line_mask_clean_valid_0 ? _GEN_852 : mask_4_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1877 = line_mask_clean_valid_0 ? _GEN_853 : mask_5_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1878 = line_mask_clean_valid_0 ? _GEN_854 : mask_6_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1879 = line_mask_clean_valid_0 ? _GEN_855 : mask_7_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1880 = line_mask_clean_valid_0 ? _GEN_856 : mask_8_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1881 = line_mask_clean_valid_0 ? _GEN_857 : mask_9_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1882 = line_mask_clean_valid_0 ? _GEN_858 : mask_10_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1883 = line_mask_clean_valid_0 ? _GEN_859 : mask_11_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1884 = line_mask_clean_valid_0 ? _GEN_860 : mask_12_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1885 = line_mask_clean_valid_0 ? _GEN_861 : mask_13_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1886 = line_mask_clean_valid_0 ? _GEN_862 : mask_14_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1887 = line_mask_clean_valid_0 ? _GEN_863 : mask_15_6_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1888 = line_mask_clean_valid_0 ? _GEN_864 : mask_0_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1889 = line_mask_clean_valid_0 ? _GEN_865 : mask_1_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1890 = line_mask_clean_valid_0 ? _GEN_866 : mask_2_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1891 = line_mask_clean_valid_0 ? _GEN_867 : mask_3_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1892 = line_mask_clean_valid_0 ? _GEN_868 : mask_4_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1893 = line_mask_clean_valid_0 ? _GEN_869 : mask_5_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1894 = line_mask_clean_valid_0 ? _GEN_870 : mask_6_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1895 = line_mask_clean_valid_0 ? _GEN_871 : mask_7_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1896 = line_mask_clean_valid_0 ? _GEN_872 : mask_8_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1897 = line_mask_clean_valid_0 ? _GEN_873 : mask_9_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1898 = line_mask_clean_valid_0 ? _GEN_874 : mask_10_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1899 = line_mask_clean_valid_0 ? _GEN_875 : mask_11_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1900 = line_mask_clean_valid_0 ? _GEN_876 : mask_12_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1901 = line_mask_clean_valid_0 ? _GEN_877 : mask_13_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1902 = line_mask_clean_valid_0 ? _GEN_878 : mask_14_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1903 = line_mask_clean_valid_0 ? _GEN_879 : mask_15_6_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1904 = line_mask_clean_valid_0 ? _GEN_880 : mask_0_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1905 = line_mask_clean_valid_0 ? _GEN_881 : mask_1_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1906 = line_mask_clean_valid_0 ? _GEN_882 : mask_2_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1907 = line_mask_clean_valid_0 ? _GEN_883 : mask_3_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1908 = line_mask_clean_valid_0 ? _GEN_884 : mask_4_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1909 = line_mask_clean_valid_0 ? _GEN_885 : mask_5_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1910 = line_mask_clean_valid_0 ? _GEN_886 : mask_6_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1911 = line_mask_clean_valid_0 ? _GEN_887 : mask_7_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1912 = line_mask_clean_valid_0 ? _GEN_888 : mask_8_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1913 = line_mask_clean_valid_0 ? _GEN_889 : mask_9_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1914 = line_mask_clean_valid_0 ? _GEN_890 : mask_10_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1915 = line_mask_clean_valid_0 ? _GEN_891 : mask_11_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1916 = line_mask_clean_valid_0 ? _GEN_892 : mask_12_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1917 = line_mask_clean_valid_0 ? _GEN_893 : mask_13_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1918 = line_mask_clean_valid_0 ? _GEN_894 : mask_14_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1919 = line_mask_clean_valid_0 ? _GEN_895 : mask_15_6_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1920 = line_mask_clean_valid_0 ? _GEN_896 : mask_0_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1921 = line_mask_clean_valid_0 ? _GEN_897 : mask_1_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1922 = line_mask_clean_valid_0 ? _GEN_898 : mask_2_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1923 = line_mask_clean_valid_0 ? _GEN_899 : mask_3_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1924 = line_mask_clean_valid_0 ? _GEN_900 : mask_4_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1925 = line_mask_clean_valid_0 ? _GEN_901 : mask_5_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1926 = line_mask_clean_valid_0 ? _GEN_902 : mask_6_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1927 = line_mask_clean_valid_0 ? _GEN_903 : mask_7_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1928 = line_mask_clean_valid_0 ? _GEN_904 : mask_8_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1929 = line_mask_clean_valid_0 ? _GEN_905 : mask_9_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1930 = line_mask_clean_valid_0 ? _GEN_906 : mask_10_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1931 = line_mask_clean_valid_0 ? _GEN_907 : mask_11_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1932 = line_mask_clean_valid_0 ? _GEN_908 : mask_12_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1933 = line_mask_clean_valid_0 ? _GEN_909 : mask_13_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1934 = line_mask_clean_valid_0 ? _GEN_910 : mask_14_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1935 = line_mask_clean_valid_0 ? _GEN_911 : mask_15_7_0; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1936 = line_mask_clean_valid_0 ? _GEN_912 : mask_0_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1937 = line_mask_clean_valid_0 ? _GEN_913 : mask_1_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1938 = line_mask_clean_valid_0 ? _GEN_914 : mask_2_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1939 = line_mask_clean_valid_0 ? _GEN_915 : mask_3_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1940 = line_mask_clean_valid_0 ? _GEN_916 : mask_4_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1941 = line_mask_clean_valid_0 ? _GEN_917 : mask_5_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1942 = line_mask_clean_valid_0 ? _GEN_918 : mask_6_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1943 = line_mask_clean_valid_0 ? _GEN_919 : mask_7_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1944 = line_mask_clean_valid_0 ? _GEN_920 : mask_8_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1945 = line_mask_clean_valid_0 ? _GEN_921 : mask_9_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1946 = line_mask_clean_valid_0 ? _GEN_922 : mask_10_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1947 = line_mask_clean_valid_0 ? _GEN_923 : mask_11_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1948 = line_mask_clean_valid_0 ? _GEN_924 : mask_12_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1949 = line_mask_clean_valid_0 ? _GEN_925 : mask_13_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1950 = line_mask_clean_valid_0 ? _GEN_926 : mask_14_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1951 = line_mask_clean_valid_0 ? _GEN_927 : mask_15_7_1; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1952 = line_mask_clean_valid_0 ? _GEN_928 : mask_0_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1953 = line_mask_clean_valid_0 ? _GEN_929 : mask_1_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1954 = line_mask_clean_valid_0 ? _GEN_930 : mask_2_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1955 = line_mask_clean_valid_0 ? _GEN_931 : mask_3_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1956 = line_mask_clean_valid_0 ? _GEN_932 : mask_4_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1957 = line_mask_clean_valid_0 ? _GEN_933 : mask_5_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1958 = line_mask_clean_valid_0 ? _GEN_934 : mask_6_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1959 = line_mask_clean_valid_0 ? _GEN_935 : mask_7_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1960 = line_mask_clean_valid_0 ? _GEN_936 : mask_8_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1961 = line_mask_clean_valid_0 ? _GEN_937 : mask_9_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1962 = line_mask_clean_valid_0 ? _GEN_938 : mask_10_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1963 = line_mask_clean_valid_0 ? _GEN_939 : mask_11_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1964 = line_mask_clean_valid_0 ? _GEN_940 : mask_12_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1965 = line_mask_clean_valid_0 ? _GEN_941 : mask_13_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1966 = line_mask_clean_valid_0 ? _GEN_942 : mask_14_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1967 = line_mask_clean_valid_0 ? _GEN_943 : mask_15_7_2; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1968 = line_mask_clean_valid_0 ? _GEN_944 : mask_0_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1969 = line_mask_clean_valid_0 ? _GEN_945 : mask_1_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1970 = line_mask_clean_valid_0 ? _GEN_946 : mask_2_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1971 = line_mask_clean_valid_0 ? _GEN_947 : mask_3_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1972 = line_mask_clean_valid_0 ? _GEN_948 : mask_4_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1973 = line_mask_clean_valid_0 ? _GEN_949 : mask_5_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1974 = line_mask_clean_valid_0 ? _GEN_950 : mask_6_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1975 = line_mask_clean_valid_0 ? _GEN_951 : mask_7_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1976 = line_mask_clean_valid_0 ? _GEN_952 : mask_8_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1977 = line_mask_clean_valid_0 ? _GEN_953 : mask_9_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1978 = line_mask_clean_valid_0 ? _GEN_954 : mask_10_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1979 = line_mask_clean_valid_0 ? _GEN_955 : mask_11_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1980 = line_mask_clean_valid_0 ? _GEN_956 : mask_12_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1981 = line_mask_clean_valid_0 ? _GEN_957 : mask_13_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1982 = line_mask_clean_valid_0 ? _GEN_958 : mask_14_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1983 = line_mask_clean_valid_0 ? _GEN_959 : mask_15_7_3; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1984 = line_mask_clean_valid_0 ? _GEN_960 : mask_0_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1985 = line_mask_clean_valid_0 ? _GEN_961 : mask_1_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1986 = line_mask_clean_valid_0 ? _GEN_962 : mask_2_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1987 = line_mask_clean_valid_0 ? _GEN_963 : mask_3_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1988 = line_mask_clean_valid_0 ? _GEN_964 : mask_4_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1989 = line_mask_clean_valid_0 ? _GEN_965 : mask_5_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1990 = line_mask_clean_valid_0 ? _GEN_966 : mask_6_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1991 = line_mask_clean_valid_0 ? _GEN_967 : mask_7_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1992 = line_mask_clean_valid_0 ? _GEN_968 : mask_8_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1993 = line_mask_clean_valid_0 ? _GEN_969 : mask_9_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1994 = line_mask_clean_valid_0 ? _GEN_970 : mask_10_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1995 = line_mask_clean_valid_0 ? _GEN_971 : mask_11_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1996 = line_mask_clean_valid_0 ? _GEN_972 : mask_12_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1997 = line_mask_clean_valid_0 ? _GEN_973 : mask_13_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1998 = line_mask_clean_valid_0 ? _GEN_974 : mask_14_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_1999 = line_mask_clean_valid_0 ? _GEN_975 : mask_15_7_4; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2000 = line_mask_clean_valid_0 ? _GEN_976 : mask_0_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2001 = line_mask_clean_valid_0 ? _GEN_977 : mask_1_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2002 = line_mask_clean_valid_0 ? _GEN_978 : mask_2_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2003 = line_mask_clean_valid_0 ? _GEN_979 : mask_3_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2004 = line_mask_clean_valid_0 ? _GEN_980 : mask_4_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2005 = line_mask_clean_valid_0 ? _GEN_981 : mask_5_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2006 = line_mask_clean_valid_0 ? _GEN_982 : mask_6_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2007 = line_mask_clean_valid_0 ? _GEN_983 : mask_7_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2008 = line_mask_clean_valid_0 ? _GEN_984 : mask_8_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2009 = line_mask_clean_valid_0 ? _GEN_985 : mask_9_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2010 = line_mask_clean_valid_0 ? _GEN_986 : mask_10_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2011 = line_mask_clean_valid_0 ? _GEN_987 : mask_11_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2012 = line_mask_clean_valid_0 ? _GEN_988 : mask_12_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2013 = line_mask_clean_valid_0 ? _GEN_989 : mask_13_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2014 = line_mask_clean_valid_0 ? _GEN_990 : mask_14_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2015 = line_mask_clean_valid_0 ? _GEN_991 : mask_15_7_5; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2016 = line_mask_clean_valid_0 ? _GEN_992 : mask_0_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2017 = line_mask_clean_valid_0 ? _GEN_993 : mask_1_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2018 = line_mask_clean_valid_0 ? _GEN_994 : mask_2_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2019 = line_mask_clean_valid_0 ? _GEN_995 : mask_3_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2020 = line_mask_clean_valid_0 ? _GEN_996 : mask_4_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2021 = line_mask_clean_valid_0 ? _GEN_997 : mask_5_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2022 = line_mask_clean_valid_0 ? _GEN_998 : mask_6_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2023 = line_mask_clean_valid_0 ? _GEN_999 : mask_7_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2024 = line_mask_clean_valid_0 ? _GEN_1000 : mask_8_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2025 = line_mask_clean_valid_0 ? _GEN_1001 : mask_9_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2026 = line_mask_clean_valid_0 ? _GEN_1002 : mask_10_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2027 = line_mask_clean_valid_0 ? _GEN_1003 : mask_11_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2028 = line_mask_clean_valid_0 ? _GEN_1004 : mask_12_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2029 = line_mask_clean_valid_0 ? _GEN_1005 : mask_13_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2030 = line_mask_clean_valid_0 ? _GEN_1006 : mask_14_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2031 = line_mask_clean_valid_0 ? _GEN_1007 : mask_15_7_6; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2032 = line_mask_clean_valid_0 ? _GEN_1008 : mask_0_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2033 = line_mask_clean_valid_0 ? _GEN_1009 : mask_1_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2034 = line_mask_clean_valid_0 ? _GEN_1010 : mask_2_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2035 = line_mask_clean_valid_0 ? _GEN_1011 : mask_3_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2036 = line_mask_clean_valid_0 ? _GEN_1012 : mask_4_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2037 = line_mask_clean_valid_0 ? _GEN_1013 : mask_5_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2038 = line_mask_clean_valid_0 ? _GEN_1014 : mask_6_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2039 = line_mask_clean_valid_0 ? _GEN_1015 : mask_7_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2040 = line_mask_clean_valid_0 ? _GEN_1016 : mask_8_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2041 = line_mask_clean_valid_0 ? _GEN_1017 : mask_9_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2042 = line_mask_clean_valid_0 ? _GEN_1018 : mask_10_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2043 = line_mask_clean_valid_0 ? _GEN_1019 : mask_11_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2044 = line_mask_clean_valid_0 ? _GEN_1020 : mask_12_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2045 = line_mask_clean_valid_0 ? _GEN_1021 : mask_13_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2046 = line_mask_clean_valid_0 ? _GEN_1022 : mask_14_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2047 = line_mask_clean_valid_0 ? _GEN_1023 : mask_15_7_7; // @[Sbuffer.scala 134:17 98:21]
  wire  _GEN_2048 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1024; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2049 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1025; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2050 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1026; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2051 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1027; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2052 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1028; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2053 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1029; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2054 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1030; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2055 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1031; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2056 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1032; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2057 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1033; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2058 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1034; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2059 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1035; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2060 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1036; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2061 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1037; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2062 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1038; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2063 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1039; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2064 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1040; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2065 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1041; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2066 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1042; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2067 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1043; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2068 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1044; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2069 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1045; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2070 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1046; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2071 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1047; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2072 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1048; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2073 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1049; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2074 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1050; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2075 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1051; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2076 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1052; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2077 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1053; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2078 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1054; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2079 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1055; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2080 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1056; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2081 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1057; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2082 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1058; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2083 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1059; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2084 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1060; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2085 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1061; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2086 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1062; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2087 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1063; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2088 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1064; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2089 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1065; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2090 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1066; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2091 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1067; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2092 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1068; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2093 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1069; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2094 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1070; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2095 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1071; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2096 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1072; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2097 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1073; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2098 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1074; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2099 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1075; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2100 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1076; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2101 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1077; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2102 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1078; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2103 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1079; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2104 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1080; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2105 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1081; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2106 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1082; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2107 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1083; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2108 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1084; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2109 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1085; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2110 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1086; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2111 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1087; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2112 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1088; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2113 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1089; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2114 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1090; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2115 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1091; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2116 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1092; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2117 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1093; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2118 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1094; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2119 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1095; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2120 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1096; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2121 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1097; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2122 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1098; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2123 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1099; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2124 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1100; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2125 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1101; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2126 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1102; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2127 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1103; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2128 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1104; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2129 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1105; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2130 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1106; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2131 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1107; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2132 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1108; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2133 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1109; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2134 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1110; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2135 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1111; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2136 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1112; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2137 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1113; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2138 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1114; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2139 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1115; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2140 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1116; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2141 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1117; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2142 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1118; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2143 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1119; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2144 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1120; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2145 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1121; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2146 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1122; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2147 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1123; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2148 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1124; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2149 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1125; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2150 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1126; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2151 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1127; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2152 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1128; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2153 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1129; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2154 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1130; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2155 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1131; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2156 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1132; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2157 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1133; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2158 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1134; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2159 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1135; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2160 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1136; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2161 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1137; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2162 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1138; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2163 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1139; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2164 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1140; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2165 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1141; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2166 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1142; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2167 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1143; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2168 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1144; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2169 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1145; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2170 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1146; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2171 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1147; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2172 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1148; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2173 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1149; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2174 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1150; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2175 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1151; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2176 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1152; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2177 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1153; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2178 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1154; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2179 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1155; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2180 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1156; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2181 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1157; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2182 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1158; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2183 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1159; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2184 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1160; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2185 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1161; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2186 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1162; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2187 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1163; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2188 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1164; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2189 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1165; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2190 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1166; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2191 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1167; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2192 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1168; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2193 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1169; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2194 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1170; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2195 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1171; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2196 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1172; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2197 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1173; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2198 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1174; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2199 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1175; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2200 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1176; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2201 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1177; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2202 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1178; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2203 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1179; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2204 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1180; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2205 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1181; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2206 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1182; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2207 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1183; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2208 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1184; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2209 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1185; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2210 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1186; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2211 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1187; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2212 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1188; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2213 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1189; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2214 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1190; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2215 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1191; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2216 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1192; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2217 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1193; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2218 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1194; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2219 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1195; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2220 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1196; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2221 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1197; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2222 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1198; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2223 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1199; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2224 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1200; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2225 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1201; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2226 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1202; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2227 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1203; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2228 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1204; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2229 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1205; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2230 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1206; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2231 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1207; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2232 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1208; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2233 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1209; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2234 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1210; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2235 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1211; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2236 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1212; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2237 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1213; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2238 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1214; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2239 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1215; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2240 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1216; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2241 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1217; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2242 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1218; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2243 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1219; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2244 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1220; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2245 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1221; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2246 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1222; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2247 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1223; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2248 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1224; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2249 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1225; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2250 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1226; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2251 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1227; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2252 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1228; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2253 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1229; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2254 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1230; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2255 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1231; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2256 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1232; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2257 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1233; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2258 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1234; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2259 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1235; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2260 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1236; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2261 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1237; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2262 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1238; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2263 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1239; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2264 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1240; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2265 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1241; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2266 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1242; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2267 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1243; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2268 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1244; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2269 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1245; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2270 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1246; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2271 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1247; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2272 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1248; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2273 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1249; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2274 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1250; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2275 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1251; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2276 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1252; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2277 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1253; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2278 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1254; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2279 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1255; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2280 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1256; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2281 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1257; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2282 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1258; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2283 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1259; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2284 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1260; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2285 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1261; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2286 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1262; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2287 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1263; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2288 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1264; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2289 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1265; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2290 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1266; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2291 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1267; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2292 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1268; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2293 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1269; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2294 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1270; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2295 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1271; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2296 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1272; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2297 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1273; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2298 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1274; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2299 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1275; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2300 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1276; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2301 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1277; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2302 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1278; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2303 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1279; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2304 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1280; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2305 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1281; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2306 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1282; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2307 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1283; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2308 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1284; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2309 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1285; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2310 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1286; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2311 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1287; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2312 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1288; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2313 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1289; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2314 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1290; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2315 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1291; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2316 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1292; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2317 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1293; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2318 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1294; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2319 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1295; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2320 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1296; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2321 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1297; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2322 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1298; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2323 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1299; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2324 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1300; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2325 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1301; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2326 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1302; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2327 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1303; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2328 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1304; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2329 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1305; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2330 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1306; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2331 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1307; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2332 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1308; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2333 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1309; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2334 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1310; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2335 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1311; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2336 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1312; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2337 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1313; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2338 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1314; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2339 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1315; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2340 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1316; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2341 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1317; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2342 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1318; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2343 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1319; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2344 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1320; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2345 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1321; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2346 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1322; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2347 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1323; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2348 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1324; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2349 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1325; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2350 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1326; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2351 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1327; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2352 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1328; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2353 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1329; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2354 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1330; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2355 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1331; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2356 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1332; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2357 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1333; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2358 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1334; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2359 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1335; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2360 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1336; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2361 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1337; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2362 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1338; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2363 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1339; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2364 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1340; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2365 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1341; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2366 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1342; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2367 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1343; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2368 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1344; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2369 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1345; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2370 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1346; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2371 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1347; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2372 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1348; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2373 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1349; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2374 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1350; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2375 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1351; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2376 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1352; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2377 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1353; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2378 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1354; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2379 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1355; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2380 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1356; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2381 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1357; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2382 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1358; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2383 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1359; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2384 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1360; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2385 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1361; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2386 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1362; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2387 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1363; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2388 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1364; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2389 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1365; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2390 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1366; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2391 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1367; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2392 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1368; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2393 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1369; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2394 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1370; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2395 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1371; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2396 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1372; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2397 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1373; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2398 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1374; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2399 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1375; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2400 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1376; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2401 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1377; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2402 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1378; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2403 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1379; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2404 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1380; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2405 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1381; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2406 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1382; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2407 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1383; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2408 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1384; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2409 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1385; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2410 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1386; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2411 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1387; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2412 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1388; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2413 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1389; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2414 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1390; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2415 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1391; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2416 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1392; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2417 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1393; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2418 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1394; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2419 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1395; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2420 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1396; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2421 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1397; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2422 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1398; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2423 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1399; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2424 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1400; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2425 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1401; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2426 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1402; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2427 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1403; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2428 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1404; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2429 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1405; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2430 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1406; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2431 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1407; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2432 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1408; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2433 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1409; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2434 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1410; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2435 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1411; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2436 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1412; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2437 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1413; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2438 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1414; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2439 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1415; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2440 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1416; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2441 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1417; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2442 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1418; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2443 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1419; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2444 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1420; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2445 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1421; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2446 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1422; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2447 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1423; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2448 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1424; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2449 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1425; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2450 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1426; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2451 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1427; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2452 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1428; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2453 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1429; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2454 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1430; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2455 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1431; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2456 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1432; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2457 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1433; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2458 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1434; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2459 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1435; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2460 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1436; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2461 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1437; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2462 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1438; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2463 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1439; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2464 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1440; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2465 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1441; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2466 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1442; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2467 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1443; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2468 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1444; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2469 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1445; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2470 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1446; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2471 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1447; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2472 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1448; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2473 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1449; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2474 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1450; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2475 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1451; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2476 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1452; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2477 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1453; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2478 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1454; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2479 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1455; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2480 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1456; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2481 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1457; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2482 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1458; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2483 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1459; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2484 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1460; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2485 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1461; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2486 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1462; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2487 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1463; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2488 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1464; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2489 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1465; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2490 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1466; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2491 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1467; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2492 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1468; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2493 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1469; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2494 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1470; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2495 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1471; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2496 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1472; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2497 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1473; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2498 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1474; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2499 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1475; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2500 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1476; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2501 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1477; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2502 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1478; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2503 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1479; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2504 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1480; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2505 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1481; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2506 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1482; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2507 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1483; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2508 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1484; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2509 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1485; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2510 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1486; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2511 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1487; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2512 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1488; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2513 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1489; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2514 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1490; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2515 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1491; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2516 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1492; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2517 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1493; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2518 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1494; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2519 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1495; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2520 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1496; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2521 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1497; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2522 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1498; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2523 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1499; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2524 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1500; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2525 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1501; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2526 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1502; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2527 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1503; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2528 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1504; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2529 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1505; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2530 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1506; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2531 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1507; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2532 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1508; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2533 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1509; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2534 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1510; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2535 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1511; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2536 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1512; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2537 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1513; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2538 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1514; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2539 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1515; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2540 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1516; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2541 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1517; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2542 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1518; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2543 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1519; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2544 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1520; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2545 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1521; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2546 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1522; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2547 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1523; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2548 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1524; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2549 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1525; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2550 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1526; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2551 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1527; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2552 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1528; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2553 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1529; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2554 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1530; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2555 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1531; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2556 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1532; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2557 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1533; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2558 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1534; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2559 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1535; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2560 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1536; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2561 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1537; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2562 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1538; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2563 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1539; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2564 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1540; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2565 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1541; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2566 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1542; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2567 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1543; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2568 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1544; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2569 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1545; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2570 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1546; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2571 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1547; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2572 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1548; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2573 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1549; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2574 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1550; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2575 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1551; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2576 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1552; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2577 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1553; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2578 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1554; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2579 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1555; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2580 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1556; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2581 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1557; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2582 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1558; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2583 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1559; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2584 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1560; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2585 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1561; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2586 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1562; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2587 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1563; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2588 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1564; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2589 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1565; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2590 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1566; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2591 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1567; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2592 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1568; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2593 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1569; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2594 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1570; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2595 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1571; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2596 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1572; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2597 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1573; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2598 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1574; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2599 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1575; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2600 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1576; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2601 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1577; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2602 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1578; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2603 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1579; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2604 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1580; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2605 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1581; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2606 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1582; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2607 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1583; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2608 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1584; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2609 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1585; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2610 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1586; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2611 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1587; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2612 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1588; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2613 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1589; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2614 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1590; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2615 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1591; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2616 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1592; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2617 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1593; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2618 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1594; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2619 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1595; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2620 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1596; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2621 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1597; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2622 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1598; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2623 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1599; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2624 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1600; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2625 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1601; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2626 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1602; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2627 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1603; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2628 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1604; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2629 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1605; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2630 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1606; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2631 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1607; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2632 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1608; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2633 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1609; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2634 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1610; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2635 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1611; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2636 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1612; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2637 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1613; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2638 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1614; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2639 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1615; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2640 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1616; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2641 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1617; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2642 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1618; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2643 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1619; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2644 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1620; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2645 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1621; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2646 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1622; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2647 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1623; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2648 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1624; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2649 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1625; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2650 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1626; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2651 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1627; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2652 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1628; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2653 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1629; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2654 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1630; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2655 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1631; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2656 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1632; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2657 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1633; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2658 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1634; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2659 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1635; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2660 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1636; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2661 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1637; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2662 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1638; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2663 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1639; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2664 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1640; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2665 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1641; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2666 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1642; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2667 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1643; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2668 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1644; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2669 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1645; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2670 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1646; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2671 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1647; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2672 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1648; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2673 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1649; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2674 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1650; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2675 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1651; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2676 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1652; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2677 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1653; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2678 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1654; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2679 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1655; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2680 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1656; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2681 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1657; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2682 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1658; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2683 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1659; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2684 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1660; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2685 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1661; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2686 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1662; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2687 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1663; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2688 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1664; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2689 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1665; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2690 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1666; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2691 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1667; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2692 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1668; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2693 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1669; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2694 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1670; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2695 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1671; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2696 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1672; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2697 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1673; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2698 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1674; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2699 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1675; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2700 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1676; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2701 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1677; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2702 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1678; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2703 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1679; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2704 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1680; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2705 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1681; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2706 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1682; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2707 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1683; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2708 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1684; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2709 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1685; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2710 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1686; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2711 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1687; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2712 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1688; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2713 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1689; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2714 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1690; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2715 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1691; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2716 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1692; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2717 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1693; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2718 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1694; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2719 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1695; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2720 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1696; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2721 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1697; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2722 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1698; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2723 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1699; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2724 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1700; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2725 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1701; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2726 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1702; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2727 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1703; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2728 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1704; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2729 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1705; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2730 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1706; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2731 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1707; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2732 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1708; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2733 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1709; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2734 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1710; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2735 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1711; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2736 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1712; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2737 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1713; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2738 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1714; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2739 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1715; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2740 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1716; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2741 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1717; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2742 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1718; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2743 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1719; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2744 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1720; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2745 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1721; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2746 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1722; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2747 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1723; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2748 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1724; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2749 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1725; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2750 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1726; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2751 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1727; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2752 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1728; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2753 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1729; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2754 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1730; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2755 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1731; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2756 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1732; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2757 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1733; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2758 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1734; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2759 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1735; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2760 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1736; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2761 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1737; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2762 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1738; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2763 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1739; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2764 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1740; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2765 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1741; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2766 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1742; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2767 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1743; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2768 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1744; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2769 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1745; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2770 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1746; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2771 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1747; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2772 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1748; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2773 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1749; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2774 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1750; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2775 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1751; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2776 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1752; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2777 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1753; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2778 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1754; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2779 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1755; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2780 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1756; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2781 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1757; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2782 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1758; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2783 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1759; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2784 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1760; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2785 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1761; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2786 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1762; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2787 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1763; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2788 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1764; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2789 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1765; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2790 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1766; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2791 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1767; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2792 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1768; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2793 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1769; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2794 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1770; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2795 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1771; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2796 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1772; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2797 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1773; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2798 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1774; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2799 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1775; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2800 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1776; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2801 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1777; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2802 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1778; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2803 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1779; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2804 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1780; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2805 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1781; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2806 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1782; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2807 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1783; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2808 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1784; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2809 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1785; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2810 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1786; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2811 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1787; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2812 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1788; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2813 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1789; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2814 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1790; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2815 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1791; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2816 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1792; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2817 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1793; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2818 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1794; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2819 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1795; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2820 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1796; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2821 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1797; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2822 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1798; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2823 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1799; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2824 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1800; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2825 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1801; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2826 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1802; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2827 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1803; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2828 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1804; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2829 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1805; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2830 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1806; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2831 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1807; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2832 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1808; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2833 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1809; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2834 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1810; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2835 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1811; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2836 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1812; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2837 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1813; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2838 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1814; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2839 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1815; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2840 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1816; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2841 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1817; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2842 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1818; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2843 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1819; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2844 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1820; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2845 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1821; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2846 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1822; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2847 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1823; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2848 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1824; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2849 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1825; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2850 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1826; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2851 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1827; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2852 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1828; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2853 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1829; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2854 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1830; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2855 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1831; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2856 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1832; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2857 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1833; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2858 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1834; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2859 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1835; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2860 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1836; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2861 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1837; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2862 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1838; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2863 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1839; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2864 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1840; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2865 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1841; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2866 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1842; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2867 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1843; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2868 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1844; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2869 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1845; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2870 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1846; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2871 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1847; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2872 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1848; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2873 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1849; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2874 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1850; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2875 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1851; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2876 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1852; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2877 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1853; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2878 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1854; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2879 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1855; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2880 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1856; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2881 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1857; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2882 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1858; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2883 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1859; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2884 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1860; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2885 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1861; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2886 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1862; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2887 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1863; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2888 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1864; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2889 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1865; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2890 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1866; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2891 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1867; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2892 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1868; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2893 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1869; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2894 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1870; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2895 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1871; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2896 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1872; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2897 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1873; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2898 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1874; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2899 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1875; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2900 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1876; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2901 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1877; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2902 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1878; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2903 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1879; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2904 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1880; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2905 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1881; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2906 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1882; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2907 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1883; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2908 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1884; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2909 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1885; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2910 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1886; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2911 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1887; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2912 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1888; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2913 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1889; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2914 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1890; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2915 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1891; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2916 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1892; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2917 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1893; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2918 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1894; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2919 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1895; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2920 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1896; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2921 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1897; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2922 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1898; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2923 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1899; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2924 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1900; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2925 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1901; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2926 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1902; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2927 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1903; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2928 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1904; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2929 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1905; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2930 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1906; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2931 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1907; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2932 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1908; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2933 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1909; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2934 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1910; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2935 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1911; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2936 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1912; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2937 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1913; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2938 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1914; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2939 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1915; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2940 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1916; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2941 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1917; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2942 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1918; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2943 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1919; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2944 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1920; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2945 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1921; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2946 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1922; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2947 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1923; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2948 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1924; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2949 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1925; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2950 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1926; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2951 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1927; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2952 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1928; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2953 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1929; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2954 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1930; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2955 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1931; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2956 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1932; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2957 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1933; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2958 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1934; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2959 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1935; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2960 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1936; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2961 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1937; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2962 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1938; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2963 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1939; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2964 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1940; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2965 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1941; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2966 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1942; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2967 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1943; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2968 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1944; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2969 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1945; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2970 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1946; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2971 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1947; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2972 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1948; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2973 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1949; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2974 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1950; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2975 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1951; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2976 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1952; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2977 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1953; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2978 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1954; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2979 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1955; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2980 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1956; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2981 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1957; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2982 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1958; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2983 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1959; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2984 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1960; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2985 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1961; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2986 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1962; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2987 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1963; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2988 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1964; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2989 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1965; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2990 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1966; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2991 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1967; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2992 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1968; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2993 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1969; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2994 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1970; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2995 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1971; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2996 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1972; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2997 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1973; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2998 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1974; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_2999 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1975; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3000 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1976; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3001 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1977; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3002 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1978; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3003 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1979; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3004 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1980; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3005 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1981; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3006 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1982; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3007 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1983; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3008 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_1984; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3009 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_1985; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3010 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_1986; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3011 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_1987; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3012 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_1988; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3013 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_1989; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3014 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_1990; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3015 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_1991; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3016 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_1992; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3017 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_1993; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3018 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_1994; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3019 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_1995; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3020 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_1996; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3021 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_1997; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3022 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_1998; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3023 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_1999; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3024 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_2000; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3025 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_2001; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3026 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_2002; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3027 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_2003; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3028 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_2004; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3029 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_2005; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3030 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_2006; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3031 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_2007; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3032 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_2008; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3033 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_2009; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3034 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_2010; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3035 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_2011; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3036 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_2012; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3037 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_2013; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3038 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_2014; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3039 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_2015; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3040 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_2016; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3041 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_2017; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3042 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_2018; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3043 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_2019; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3044 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_2020; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3045 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_2021; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3046 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_2022; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3047 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_2023; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3048 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_2024; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3049 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_2025; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3050 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_2026; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3051 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_2027; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3052 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_2028; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3053 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_2029; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3054 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_2030; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3055 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_2031; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3056 = 4'h0 == line_mask_clean_line_1 ? 1'h0 : _GEN_2032; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3057 = 4'h1 == line_mask_clean_line_1 ? 1'h0 : _GEN_2033; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3058 = 4'h2 == line_mask_clean_line_1 ? 1'h0 : _GEN_2034; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3059 = 4'h3 == line_mask_clean_line_1 ? 1'h0 : _GEN_2035; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3060 = 4'h4 == line_mask_clean_line_1 ? 1'h0 : _GEN_2036; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3061 = 4'h5 == line_mask_clean_line_1 ? 1'h0 : _GEN_2037; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3062 = 4'h6 == line_mask_clean_line_1 ? 1'h0 : _GEN_2038; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3063 = 4'h7 == line_mask_clean_line_1 ? 1'h0 : _GEN_2039; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3064 = 4'h8 == line_mask_clean_line_1 ? 1'h0 : _GEN_2040; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3065 = 4'h9 == line_mask_clean_line_1 ? 1'h0 : _GEN_2041; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3066 = 4'ha == line_mask_clean_line_1 ? 1'h0 : _GEN_2042; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3067 = 4'hb == line_mask_clean_line_1 ? 1'h0 : _GEN_2043; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3068 = 4'hc == line_mask_clean_line_1 ? 1'h0 : _GEN_2044; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3069 = 4'hd == line_mask_clean_line_1 ? 1'h0 : _GEN_2045; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3070 = 4'he == line_mask_clean_line_1 ? 1'h0 : _GEN_2046; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3071 = 4'hf == line_mask_clean_line_1 ? 1'h0 : _GEN_2047; // @[Sbuffer.scala 137:{34,34}]
  wire  _GEN_3072 = line_mask_clean_valid_1 ? _GEN_2048 : _GEN_1024; // @[Sbuffer.scala 134:17]
  wire  _GEN_3073 = line_mask_clean_valid_1 ? _GEN_2049 : _GEN_1025; // @[Sbuffer.scala 134:17]
  wire  _GEN_3074 = line_mask_clean_valid_1 ? _GEN_2050 : _GEN_1026; // @[Sbuffer.scala 134:17]
  wire  _GEN_3075 = line_mask_clean_valid_1 ? _GEN_2051 : _GEN_1027; // @[Sbuffer.scala 134:17]
  wire  _GEN_3076 = line_mask_clean_valid_1 ? _GEN_2052 : _GEN_1028; // @[Sbuffer.scala 134:17]
  wire  _GEN_3077 = line_mask_clean_valid_1 ? _GEN_2053 : _GEN_1029; // @[Sbuffer.scala 134:17]
  wire  _GEN_3078 = line_mask_clean_valid_1 ? _GEN_2054 : _GEN_1030; // @[Sbuffer.scala 134:17]
  wire  _GEN_3079 = line_mask_clean_valid_1 ? _GEN_2055 : _GEN_1031; // @[Sbuffer.scala 134:17]
  wire  _GEN_3080 = line_mask_clean_valid_1 ? _GEN_2056 : _GEN_1032; // @[Sbuffer.scala 134:17]
  wire  _GEN_3081 = line_mask_clean_valid_1 ? _GEN_2057 : _GEN_1033; // @[Sbuffer.scala 134:17]
  wire  _GEN_3082 = line_mask_clean_valid_1 ? _GEN_2058 : _GEN_1034; // @[Sbuffer.scala 134:17]
  wire  _GEN_3083 = line_mask_clean_valid_1 ? _GEN_2059 : _GEN_1035; // @[Sbuffer.scala 134:17]
  wire  _GEN_3084 = line_mask_clean_valid_1 ? _GEN_2060 : _GEN_1036; // @[Sbuffer.scala 134:17]
  wire  _GEN_3085 = line_mask_clean_valid_1 ? _GEN_2061 : _GEN_1037; // @[Sbuffer.scala 134:17]
  wire  _GEN_3086 = line_mask_clean_valid_1 ? _GEN_2062 : _GEN_1038; // @[Sbuffer.scala 134:17]
  wire  _GEN_3087 = line_mask_clean_valid_1 ? _GEN_2063 : _GEN_1039; // @[Sbuffer.scala 134:17]
  wire  _GEN_3088 = line_mask_clean_valid_1 ? _GEN_2064 : _GEN_1040; // @[Sbuffer.scala 134:17]
  wire  _GEN_3089 = line_mask_clean_valid_1 ? _GEN_2065 : _GEN_1041; // @[Sbuffer.scala 134:17]
  wire  _GEN_3090 = line_mask_clean_valid_1 ? _GEN_2066 : _GEN_1042; // @[Sbuffer.scala 134:17]
  wire  _GEN_3091 = line_mask_clean_valid_1 ? _GEN_2067 : _GEN_1043; // @[Sbuffer.scala 134:17]
  wire  _GEN_3092 = line_mask_clean_valid_1 ? _GEN_2068 : _GEN_1044; // @[Sbuffer.scala 134:17]
  wire  _GEN_3093 = line_mask_clean_valid_1 ? _GEN_2069 : _GEN_1045; // @[Sbuffer.scala 134:17]
  wire  _GEN_3094 = line_mask_clean_valid_1 ? _GEN_2070 : _GEN_1046; // @[Sbuffer.scala 134:17]
  wire  _GEN_3095 = line_mask_clean_valid_1 ? _GEN_2071 : _GEN_1047; // @[Sbuffer.scala 134:17]
  wire  _GEN_3096 = line_mask_clean_valid_1 ? _GEN_2072 : _GEN_1048; // @[Sbuffer.scala 134:17]
  wire  _GEN_3097 = line_mask_clean_valid_1 ? _GEN_2073 : _GEN_1049; // @[Sbuffer.scala 134:17]
  wire  _GEN_3098 = line_mask_clean_valid_1 ? _GEN_2074 : _GEN_1050; // @[Sbuffer.scala 134:17]
  wire  _GEN_3099 = line_mask_clean_valid_1 ? _GEN_2075 : _GEN_1051; // @[Sbuffer.scala 134:17]
  wire  _GEN_3100 = line_mask_clean_valid_1 ? _GEN_2076 : _GEN_1052; // @[Sbuffer.scala 134:17]
  wire  _GEN_3101 = line_mask_clean_valid_1 ? _GEN_2077 : _GEN_1053; // @[Sbuffer.scala 134:17]
  wire  _GEN_3102 = line_mask_clean_valid_1 ? _GEN_2078 : _GEN_1054; // @[Sbuffer.scala 134:17]
  wire  _GEN_3103 = line_mask_clean_valid_1 ? _GEN_2079 : _GEN_1055; // @[Sbuffer.scala 134:17]
  wire  _GEN_3104 = line_mask_clean_valid_1 ? _GEN_2080 : _GEN_1056; // @[Sbuffer.scala 134:17]
  wire  _GEN_3105 = line_mask_clean_valid_1 ? _GEN_2081 : _GEN_1057; // @[Sbuffer.scala 134:17]
  wire  _GEN_3106 = line_mask_clean_valid_1 ? _GEN_2082 : _GEN_1058; // @[Sbuffer.scala 134:17]
  wire  _GEN_3107 = line_mask_clean_valid_1 ? _GEN_2083 : _GEN_1059; // @[Sbuffer.scala 134:17]
  wire  _GEN_3108 = line_mask_clean_valid_1 ? _GEN_2084 : _GEN_1060; // @[Sbuffer.scala 134:17]
  wire  _GEN_3109 = line_mask_clean_valid_1 ? _GEN_2085 : _GEN_1061; // @[Sbuffer.scala 134:17]
  wire  _GEN_3110 = line_mask_clean_valid_1 ? _GEN_2086 : _GEN_1062; // @[Sbuffer.scala 134:17]
  wire  _GEN_3111 = line_mask_clean_valid_1 ? _GEN_2087 : _GEN_1063; // @[Sbuffer.scala 134:17]
  wire  _GEN_3112 = line_mask_clean_valid_1 ? _GEN_2088 : _GEN_1064; // @[Sbuffer.scala 134:17]
  wire  _GEN_3113 = line_mask_clean_valid_1 ? _GEN_2089 : _GEN_1065; // @[Sbuffer.scala 134:17]
  wire  _GEN_3114 = line_mask_clean_valid_1 ? _GEN_2090 : _GEN_1066; // @[Sbuffer.scala 134:17]
  wire  _GEN_3115 = line_mask_clean_valid_1 ? _GEN_2091 : _GEN_1067; // @[Sbuffer.scala 134:17]
  wire  _GEN_3116 = line_mask_clean_valid_1 ? _GEN_2092 : _GEN_1068; // @[Sbuffer.scala 134:17]
  wire  _GEN_3117 = line_mask_clean_valid_1 ? _GEN_2093 : _GEN_1069; // @[Sbuffer.scala 134:17]
  wire  _GEN_3118 = line_mask_clean_valid_1 ? _GEN_2094 : _GEN_1070; // @[Sbuffer.scala 134:17]
  wire  _GEN_3119 = line_mask_clean_valid_1 ? _GEN_2095 : _GEN_1071; // @[Sbuffer.scala 134:17]
  wire  _GEN_3120 = line_mask_clean_valid_1 ? _GEN_2096 : _GEN_1072; // @[Sbuffer.scala 134:17]
  wire  _GEN_3121 = line_mask_clean_valid_1 ? _GEN_2097 : _GEN_1073; // @[Sbuffer.scala 134:17]
  wire  _GEN_3122 = line_mask_clean_valid_1 ? _GEN_2098 : _GEN_1074; // @[Sbuffer.scala 134:17]
  wire  _GEN_3123 = line_mask_clean_valid_1 ? _GEN_2099 : _GEN_1075; // @[Sbuffer.scala 134:17]
  wire  _GEN_3124 = line_mask_clean_valid_1 ? _GEN_2100 : _GEN_1076; // @[Sbuffer.scala 134:17]
  wire  _GEN_3125 = line_mask_clean_valid_1 ? _GEN_2101 : _GEN_1077; // @[Sbuffer.scala 134:17]
  wire  _GEN_3126 = line_mask_clean_valid_1 ? _GEN_2102 : _GEN_1078; // @[Sbuffer.scala 134:17]
  wire  _GEN_3127 = line_mask_clean_valid_1 ? _GEN_2103 : _GEN_1079; // @[Sbuffer.scala 134:17]
  wire  _GEN_3128 = line_mask_clean_valid_1 ? _GEN_2104 : _GEN_1080; // @[Sbuffer.scala 134:17]
  wire  _GEN_3129 = line_mask_clean_valid_1 ? _GEN_2105 : _GEN_1081; // @[Sbuffer.scala 134:17]
  wire  _GEN_3130 = line_mask_clean_valid_1 ? _GEN_2106 : _GEN_1082; // @[Sbuffer.scala 134:17]
  wire  _GEN_3131 = line_mask_clean_valid_1 ? _GEN_2107 : _GEN_1083; // @[Sbuffer.scala 134:17]
  wire  _GEN_3132 = line_mask_clean_valid_1 ? _GEN_2108 : _GEN_1084; // @[Sbuffer.scala 134:17]
  wire  _GEN_3133 = line_mask_clean_valid_1 ? _GEN_2109 : _GEN_1085; // @[Sbuffer.scala 134:17]
  wire  _GEN_3134 = line_mask_clean_valid_1 ? _GEN_2110 : _GEN_1086; // @[Sbuffer.scala 134:17]
  wire  _GEN_3135 = line_mask_clean_valid_1 ? _GEN_2111 : _GEN_1087; // @[Sbuffer.scala 134:17]
  wire  _GEN_3136 = line_mask_clean_valid_1 ? _GEN_2112 : _GEN_1088; // @[Sbuffer.scala 134:17]
  wire  _GEN_3137 = line_mask_clean_valid_1 ? _GEN_2113 : _GEN_1089; // @[Sbuffer.scala 134:17]
  wire  _GEN_3138 = line_mask_clean_valid_1 ? _GEN_2114 : _GEN_1090; // @[Sbuffer.scala 134:17]
  wire  _GEN_3139 = line_mask_clean_valid_1 ? _GEN_2115 : _GEN_1091; // @[Sbuffer.scala 134:17]
  wire  _GEN_3140 = line_mask_clean_valid_1 ? _GEN_2116 : _GEN_1092; // @[Sbuffer.scala 134:17]
  wire  _GEN_3141 = line_mask_clean_valid_1 ? _GEN_2117 : _GEN_1093; // @[Sbuffer.scala 134:17]
  wire  _GEN_3142 = line_mask_clean_valid_1 ? _GEN_2118 : _GEN_1094; // @[Sbuffer.scala 134:17]
  wire  _GEN_3143 = line_mask_clean_valid_1 ? _GEN_2119 : _GEN_1095; // @[Sbuffer.scala 134:17]
  wire  _GEN_3144 = line_mask_clean_valid_1 ? _GEN_2120 : _GEN_1096; // @[Sbuffer.scala 134:17]
  wire  _GEN_3145 = line_mask_clean_valid_1 ? _GEN_2121 : _GEN_1097; // @[Sbuffer.scala 134:17]
  wire  _GEN_3146 = line_mask_clean_valid_1 ? _GEN_2122 : _GEN_1098; // @[Sbuffer.scala 134:17]
  wire  _GEN_3147 = line_mask_clean_valid_1 ? _GEN_2123 : _GEN_1099; // @[Sbuffer.scala 134:17]
  wire  _GEN_3148 = line_mask_clean_valid_1 ? _GEN_2124 : _GEN_1100; // @[Sbuffer.scala 134:17]
  wire  _GEN_3149 = line_mask_clean_valid_1 ? _GEN_2125 : _GEN_1101; // @[Sbuffer.scala 134:17]
  wire  _GEN_3150 = line_mask_clean_valid_1 ? _GEN_2126 : _GEN_1102; // @[Sbuffer.scala 134:17]
  wire  _GEN_3151 = line_mask_clean_valid_1 ? _GEN_2127 : _GEN_1103; // @[Sbuffer.scala 134:17]
  wire  _GEN_3152 = line_mask_clean_valid_1 ? _GEN_2128 : _GEN_1104; // @[Sbuffer.scala 134:17]
  wire  _GEN_3153 = line_mask_clean_valid_1 ? _GEN_2129 : _GEN_1105; // @[Sbuffer.scala 134:17]
  wire  _GEN_3154 = line_mask_clean_valid_1 ? _GEN_2130 : _GEN_1106; // @[Sbuffer.scala 134:17]
  wire  _GEN_3155 = line_mask_clean_valid_1 ? _GEN_2131 : _GEN_1107; // @[Sbuffer.scala 134:17]
  wire  _GEN_3156 = line_mask_clean_valid_1 ? _GEN_2132 : _GEN_1108; // @[Sbuffer.scala 134:17]
  wire  _GEN_3157 = line_mask_clean_valid_1 ? _GEN_2133 : _GEN_1109; // @[Sbuffer.scala 134:17]
  wire  _GEN_3158 = line_mask_clean_valid_1 ? _GEN_2134 : _GEN_1110; // @[Sbuffer.scala 134:17]
  wire  _GEN_3159 = line_mask_clean_valid_1 ? _GEN_2135 : _GEN_1111; // @[Sbuffer.scala 134:17]
  wire  _GEN_3160 = line_mask_clean_valid_1 ? _GEN_2136 : _GEN_1112; // @[Sbuffer.scala 134:17]
  wire  _GEN_3161 = line_mask_clean_valid_1 ? _GEN_2137 : _GEN_1113; // @[Sbuffer.scala 134:17]
  wire  _GEN_3162 = line_mask_clean_valid_1 ? _GEN_2138 : _GEN_1114; // @[Sbuffer.scala 134:17]
  wire  _GEN_3163 = line_mask_clean_valid_1 ? _GEN_2139 : _GEN_1115; // @[Sbuffer.scala 134:17]
  wire  _GEN_3164 = line_mask_clean_valid_1 ? _GEN_2140 : _GEN_1116; // @[Sbuffer.scala 134:17]
  wire  _GEN_3165 = line_mask_clean_valid_1 ? _GEN_2141 : _GEN_1117; // @[Sbuffer.scala 134:17]
  wire  _GEN_3166 = line_mask_clean_valid_1 ? _GEN_2142 : _GEN_1118; // @[Sbuffer.scala 134:17]
  wire  _GEN_3167 = line_mask_clean_valid_1 ? _GEN_2143 : _GEN_1119; // @[Sbuffer.scala 134:17]
  wire  _GEN_3168 = line_mask_clean_valid_1 ? _GEN_2144 : _GEN_1120; // @[Sbuffer.scala 134:17]
  wire  _GEN_3169 = line_mask_clean_valid_1 ? _GEN_2145 : _GEN_1121; // @[Sbuffer.scala 134:17]
  wire  _GEN_3170 = line_mask_clean_valid_1 ? _GEN_2146 : _GEN_1122; // @[Sbuffer.scala 134:17]
  wire  _GEN_3171 = line_mask_clean_valid_1 ? _GEN_2147 : _GEN_1123; // @[Sbuffer.scala 134:17]
  wire  _GEN_3172 = line_mask_clean_valid_1 ? _GEN_2148 : _GEN_1124; // @[Sbuffer.scala 134:17]
  wire  _GEN_3173 = line_mask_clean_valid_1 ? _GEN_2149 : _GEN_1125; // @[Sbuffer.scala 134:17]
  wire  _GEN_3174 = line_mask_clean_valid_1 ? _GEN_2150 : _GEN_1126; // @[Sbuffer.scala 134:17]
  wire  _GEN_3175 = line_mask_clean_valid_1 ? _GEN_2151 : _GEN_1127; // @[Sbuffer.scala 134:17]
  wire  _GEN_3176 = line_mask_clean_valid_1 ? _GEN_2152 : _GEN_1128; // @[Sbuffer.scala 134:17]
  wire  _GEN_3177 = line_mask_clean_valid_1 ? _GEN_2153 : _GEN_1129; // @[Sbuffer.scala 134:17]
  wire  _GEN_3178 = line_mask_clean_valid_1 ? _GEN_2154 : _GEN_1130; // @[Sbuffer.scala 134:17]
  wire  _GEN_3179 = line_mask_clean_valid_1 ? _GEN_2155 : _GEN_1131; // @[Sbuffer.scala 134:17]
  wire  _GEN_3180 = line_mask_clean_valid_1 ? _GEN_2156 : _GEN_1132; // @[Sbuffer.scala 134:17]
  wire  _GEN_3181 = line_mask_clean_valid_1 ? _GEN_2157 : _GEN_1133; // @[Sbuffer.scala 134:17]
  wire  _GEN_3182 = line_mask_clean_valid_1 ? _GEN_2158 : _GEN_1134; // @[Sbuffer.scala 134:17]
  wire  _GEN_3183 = line_mask_clean_valid_1 ? _GEN_2159 : _GEN_1135; // @[Sbuffer.scala 134:17]
  wire  _GEN_3184 = line_mask_clean_valid_1 ? _GEN_2160 : _GEN_1136; // @[Sbuffer.scala 134:17]
  wire  _GEN_3185 = line_mask_clean_valid_1 ? _GEN_2161 : _GEN_1137; // @[Sbuffer.scala 134:17]
  wire  _GEN_3186 = line_mask_clean_valid_1 ? _GEN_2162 : _GEN_1138; // @[Sbuffer.scala 134:17]
  wire  _GEN_3187 = line_mask_clean_valid_1 ? _GEN_2163 : _GEN_1139; // @[Sbuffer.scala 134:17]
  wire  _GEN_3188 = line_mask_clean_valid_1 ? _GEN_2164 : _GEN_1140; // @[Sbuffer.scala 134:17]
  wire  _GEN_3189 = line_mask_clean_valid_1 ? _GEN_2165 : _GEN_1141; // @[Sbuffer.scala 134:17]
  wire  _GEN_3190 = line_mask_clean_valid_1 ? _GEN_2166 : _GEN_1142; // @[Sbuffer.scala 134:17]
  wire  _GEN_3191 = line_mask_clean_valid_1 ? _GEN_2167 : _GEN_1143; // @[Sbuffer.scala 134:17]
  wire  _GEN_3192 = line_mask_clean_valid_1 ? _GEN_2168 : _GEN_1144; // @[Sbuffer.scala 134:17]
  wire  _GEN_3193 = line_mask_clean_valid_1 ? _GEN_2169 : _GEN_1145; // @[Sbuffer.scala 134:17]
  wire  _GEN_3194 = line_mask_clean_valid_1 ? _GEN_2170 : _GEN_1146; // @[Sbuffer.scala 134:17]
  wire  _GEN_3195 = line_mask_clean_valid_1 ? _GEN_2171 : _GEN_1147; // @[Sbuffer.scala 134:17]
  wire  _GEN_3196 = line_mask_clean_valid_1 ? _GEN_2172 : _GEN_1148; // @[Sbuffer.scala 134:17]
  wire  _GEN_3197 = line_mask_clean_valid_1 ? _GEN_2173 : _GEN_1149; // @[Sbuffer.scala 134:17]
  wire  _GEN_3198 = line_mask_clean_valid_1 ? _GEN_2174 : _GEN_1150; // @[Sbuffer.scala 134:17]
  wire  _GEN_3199 = line_mask_clean_valid_1 ? _GEN_2175 : _GEN_1151; // @[Sbuffer.scala 134:17]
  wire  _GEN_3200 = line_mask_clean_valid_1 ? _GEN_2176 : _GEN_1152; // @[Sbuffer.scala 134:17]
  wire  _GEN_3201 = line_mask_clean_valid_1 ? _GEN_2177 : _GEN_1153; // @[Sbuffer.scala 134:17]
  wire  _GEN_3202 = line_mask_clean_valid_1 ? _GEN_2178 : _GEN_1154; // @[Sbuffer.scala 134:17]
  wire  _GEN_3203 = line_mask_clean_valid_1 ? _GEN_2179 : _GEN_1155; // @[Sbuffer.scala 134:17]
  wire  _GEN_3204 = line_mask_clean_valid_1 ? _GEN_2180 : _GEN_1156; // @[Sbuffer.scala 134:17]
  wire  _GEN_3205 = line_mask_clean_valid_1 ? _GEN_2181 : _GEN_1157; // @[Sbuffer.scala 134:17]
  wire  _GEN_3206 = line_mask_clean_valid_1 ? _GEN_2182 : _GEN_1158; // @[Sbuffer.scala 134:17]
  wire  _GEN_3207 = line_mask_clean_valid_1 ? _GEN_2183 : _GEN_1159; // @[Sbuffer.scala 134:17]
  wire  _GEN_3208 = line_mask_clean_valid_1 ? _GEN_2184 : _GEN_1160; // @[Sbuffer.scala 134:17]
  wire  _GEN_3209 = line_mask_clean_valid_1 ? _GEN_2185 : _GEN_1161; // @[Sbuffer.scala 134:17]
  wire  _GEN_3210 = line_mask_clean_valid_1 ? _GEN_2186 : _GEN_1162; // @[Sbuffer.scala 134:17]
  wire  _GEN_3211 = line_mask_clean_valid_1 ? _GEN_2187 : _GEN_1163; // @[Sbuffer.scala 134:17]
  wire  _GEN_3212 = line_mask_clean_valid_1 ? _GEN_2188 : _GEN_1164; // @[Sbuffer.scala 134:17]
  wire  _GEN_3213 = line_mask_clean_valid_1 ? _GEN_2189 : _GEN_1165; // @[Sbuffer.scala 134:17]
  wire  _GEN_3214 = line_mask_clean_valid_1 ? _GEN_2190 : _GEN_1166; // @[Sbuffer.scala 134:17]
  wire  _GEN_3215 = line_mask_clean_valid_1 ? _GEN_2191 : _GEN_1167; // @[Sbuffer.scala 134:17]
  wire  _GEN_3216 = line_mask_clean_valid_1 ? _GEN_2192 : _GEN_1168; // @[Sbuffer.scala 134:17]
  wire  _GEN_3217 = line_mask_clean_valid_1 ? _GEN_2193 : _GEN_1169; // @[Sbuffer.scala 134:17]
  wire  _GEN_3218 = line_mask_clean_valid_1 ? _GEN_2194 : _GEN_1170; // @[Sbuffer.scala 134:17]
  wire  _GEN_3219 = line_mask_clean_valid_1 ? _GEN_2195 : _GEN_1171; // @[Sbuffer.scala 134:17]
  wire  _GEN_3220 = line_mask_clean_valid_1 ? _GEN_2196 : _GEN_1172; // @[Sbuffer.scala 134:17]
  wire  _GEN_3221 = line_mask_clean_valid_1 ? _GEN_2197 : _GEN_1173; // @[Sbuffer.scala 134:17]
  wire  _GEN_3222 = line_mask_clean_valid_1 ? _GEN_2198 : _GEN_1174; // @[Sbuffer.scala 134:17]
  wire  _GEN_3223 = line_mask_clean_valid_1 ? _GEN_2199 : _GEN_1175; // @[Sbuffer.scala 134:17]
  wire  _GEN_3224 = line_mask_clean_valid_1 ? _GEN_2200 : _GEN_1176; // @[Sbuffer.scala 134:17]
  wire  _GEN_3225 = line_mask_clean_valid_1 ? _GEN_2201 : _GEN_1177; // @[Sbuffer.scala 134:17]
  wire  _GEN_3226 = line_mask_clean_valid_1 ? _GEN_2202 : _GEN_1178; // @[Sbuffer.scala 134:17]
  wire  _GEN_3227 = line_mask_clean_valid_1 ? _GEN_2203 : _GEN_1179; // @[Sbuffer.scala 134:17]
  wire  _GEN_3228 = line_mask_clean_valid_1 ? _GEN_2204 : _GEN_1180; // @[Sbuffer.scala 134:17]
  wire  _GEN_3229 = line_mask_clean_valid_1 ? _GEN_2205 : _GEN_1181; // @[Sbuffer.scala 134:17]
  wire  _GEN_3230 = line_mask_clean_valid_1 ? _GEN_2206 : _GEN_1182; // @[Sbuffer.scala 134:17]
  wire  _GEN_3231 = line_mask_clean_valid_1 ? _GEN_2207 : _GEN_1183; // @[Sbuffer.scala 134:17]
  wire  _GEN_3232 = line_mask_clean_valid_1 ? _GEN_2208 : _GEN_1184; // @[Sbuffer.scala 134:17]
  wire  _GEN_3233 = line_mask_clean_valid_1 ? _GEN_2209 : _GEN_1185; // @[Sbuffer.scala 134:17]
  wire  _GEN_3234 = line_mask_clean_valid_1 ? _GEN_2210 : _GEN_1186; // @[Sbuffer.scala 134:17]
  wire  _GEN_3235 = line_mask_clean_valid_1 ? _GEN_2211 : _GEN_1187; // @[Sbuffer.scala 134:17]
  wire  _GEN_3236 = line_mask_clean_valid_1 ? _GEN_2212 : _GEN_1188; // @[Sbuffer.scala 134:17]
  wire  _GEN_3237 = line_mask_clean_valid_1 ? _GEN_2213 : _GEN_1189; // @[Sbuffer.scala 134:17]
  wire  _GEN_3238 = line_mask_clean_valid_1 ? _GEN_2214 : _GEN_1190; // @[Sbuffer.scala 134:17]
  wire  _GEN_3239 = line_mask_clean_valid_1 ? _GEN_2215 : _GEN_1191; // @[Sbuffer.scala 134:17]
  wire  _GEN_3240 = line_mask_clean_valid_1 ? _GEN_2216 : _GEN_1192; // @[Sbuffer.scala 134:17]
  wire  _GEN_3241 = line_mask_clean_valid_1 ? _GEN_2217 : _GEN_1193; // @[Sbuffer.scala 134:17]
  wire  _GEN_3242 = line_mask_clean_valid_1 ? _GEN_2218 : _GEN_1194; // @[Sbuffer.scala 134:17]
  wire  _GEN_3243 = line_mask_clean_valid_1 ? _GEN_2219 : _GEN_1195; // @[Sbuffer.scala 134:17]
  wire  _GEN_3244 = line_mask_clean_valid_1 ? _GEN_2220 : _GEN_1196; // @[Sbuffer.scala 134:17]
  wire  _GEN_3245 = line_mask_clean_valid_1 ? _GEN_2221 : _GEN_1197; // @[Sbuffer.scala 134:17]
  wire  _GEN_3246 = line_mask_clean_valid_1 ? _GEN_2222 : _GEN_1198; // @[Sbuffer.scala 134:17]
  wire  _GEN_3247 = line_mask_clean_valid_1 ? _GEN_2223 : _GEN_1199; // @[Sbuffer.scala 134:17]
  wire  _GEN_3248 = line_mask_clean_valid_1 ? _GEN_2224 : _GEN_1200; // @[Sbuffer.scala 134:17]
  wire  _GEN_3249 = line_mask_clean_valid_1 ? _GEN_2225 : _GEN_1201; // @[Sbuffer.scala 134:17]
  wire  _GEN_3250 = line_mask_clean_valid_1 ? _GEN_2226 : _GEN_1202; // @[Sbuffer.scala 134:17]
  wire  _GEN_3251 = line_mask_clean_valid_1 ? _GEN_2227 : _GEN_1203; // @[Sbuffer.scala 134:17]
  wire  _GEN_3252 = line_mask_clean_valid_1 ? _GEN_2228 : _GEN_1204; // @[Sbuffer.scala 134:17]
  wire  _GEN_3253 = line_mask_clean_valid_1 ? _GEN_2229 : _GEN_1205; // @[Sbuffer.scala 134:17]
  wire  _GEN_3254 = line_mask_clean_valid_1 ? _GEN_2230 : _GEN_1206; // @[Sbuffer.scala 134:17]
  wire  _GEN_3255 = line_mask_clean_valid_1 ? _GEN_2231 : _GEN_1207; // @[Sbuffer.scala 134:17]
  wire  _GEN_3256 = line_mask_clean_valid_1 ? _GEN_2232 : _GEN_1208; // @[Sbuffer.scala 134:17]
  wire  _GEN_3257 = line_mask_clean_valid_1 ? _GEN_2233 : _GEN_1209; // @[Sbuffer.scala 134:17]
  wire  _GEN_3258 = line_mask_clean_valid_1 ? _GEN_2234 : _GEN_1210; // @[Sbuffer.scala 134:17]
  wire  _GEN_3259 = line_mask_clean_valid_1 ? _GEN_2235 : _GEN_1211; // @[Sbuffer.scala 134:17]
  wire  _GEN_3260 = line_mask_clean_valid_1 ? _GEN_2236 : _GEN_1212; // @[Sbuffer.scala 134:17]
  wire  _GEN_3261 = line_mask_clean_valid_1 ? _GEN_2237 : _GEN_1213; // @[Sbuffer.scala 134:17]
  wire  _GEN_3262 = line_mask_clean_valid_1 ? _GEN_2238 : _GEN_1214; // @[Sbuffer.scala 134:17]
  wire  _GEN_3263 = line_mask_clean_valid_1 ? _GEN_2239 : _GEN_1215; // @[Sbuffer.scala 134:17]
  wire  _GEN_3264 = line_mask_clean_valid_1 ? _GEN_2240 : _GEN_1216; // @[Sbuffer.scala 134:17]
  wire  _GEN_3265 = line_mask_clean_valid_1 ? _GEN_2241 : _GEN_1217; // @[Sbuffer.scala 134:17]
  wire  _GEN_3266 = line_mask_clean_valid_1 ? _GEN_2242 : _GEN_1218; // @[Sbuffer.scala 134:17]
  wire  _GEN_3267 = line_mask_clean_valid_1 ? _GEN_2243 : _GEN_1219; // @[Sbuffer.scala 134:17]
  wire  _GEN_3268 = line_mask_clean_valid_1 ? _GEN_2244 : _GEN_1220; // @[Sbuffer.scala 134:17]
  wire  _GEN_3269 = line_mask_clean_valid_1 ? _GEN_2245 : _GEN_1221; // @[Sbuffer.scala 134:17]
  wire  _GEN_3270 = line_mask_clean_valid_1 ? _GEN_2246 : _GEN_1222; // @[Sbuffer.scala 134:17]
  wire  _GEN_3271 = line_mask_clean_valid_1 ? _GEN_2247 : _GEN_1223; // @[Sbuffer.scala 134:17]
  wire  _GEN_3272 = line_mask_clean_valid_1 ? _GEN_2248 : _GEN_1224; // @[Sbuffer.scala 134:17]
  wire  _GEN_3273 = line_mask_clean_valid_1 ? _GEN_2249 : _GEN_1225; // @[Sbuffer.scala 134:17]
  wire  _GEN_3274 = line_mask_clean_valid_1 ? _GEN_2250 : _GEN_1226; // @[Sbuffer.scala 134:17]
  wire  _GEN_3275 = line_mask_clean_valid_1 ? _GEN_2251 : _GEN_1227; // @[Sbuffer.scala 134:17]
  wire  _GEN_3276 = line_mask_clean_valid_1 ? _GEN_2252 : _GEN_1228; // @[Sbuffer.scala 134:17]
  wire  _GEN_3277 = line_mask_clean_valid_1 ? _GEN_2253 : _GEN_1229; // @[Sbuffer.scala 134:17]
  wire  _GEN_3278 = line_mask_clean_valid_1 ? _GEN_2254 : _GEN_1230; // @[Sbuffer.scala 134:17]
  wire  _GEN_3279 = line_mask_clean_valid_1 ? _GEN_2255 : _GEN_1231; // @[Sbuffer.scala 134:17]
  wire  _GEN_3280 = line_mask_clean_valid_1 ? _GEN_2256 : _GEN_1232; // @[Sbuffer.scala 134:17]
  wire  _GEN_3281 = line_mask_clean_valid_1 ? _GEN_2257 : _GEN_1233; // @[Sbuffer.scala 134:17]
  wire  _GEN_3282 = line_mask_clean_valid_1 ? _GEN_2258 : _GEN_1234; // @[Sbuffer.scala 134:17]
  wire  _GEN_3283 = line_mask_clean_valid_1 ? _GEN_2259 : _GEN_1235; // @[Sbuffer.scala 134:17]
  wire  _GEN_3284 = line_mask_clean_valid_1 ? _GEN_2260 : _GEN_1236; // @[Sbuffer.scala 134:17]
  wire  _GEN_3285 = line_mask_clean_valid_1 ? _GEN_2261 : _GEN_1237; // @[Sbuffer.scala 134:17]
  wire  _GEN_3286 = line_mask_clean_valid_1 ? _GEN_2262 : _GEN_1238; // @[Sbuffer.scala 134:17]
  wire  _GEN_3287 = line_mask_clean_valid_1 ? _GEN_2263 : _GEN_1239; // @[Sbuffer.scala 134:17]
  wire  _GEN_3288 = line_mask_clean_valid_1 ? _GEN_2264 : _GEN_1240; // @[Sbuffer.scala 134:17]
  wire  _GEN_3289 = line_mask_clean_valid_1 ? _GEN_2265 : _GEN_1241; // @[Sbuffer.scala 134:17]
  wire  _GEN_3290 = line_mask_clean_valid_1 ? _GEN_2266 : _GEN_1242; // @[Sbuffer.scala 134:17]
  wire  _GEN_3291 = line_mask_clean_valid_1 ? _GEN_2267 : _GEN_1243; // @[Sbuffer.scala 134:17]
  wire  _GEN_3292 = line_mask_clean_valid_1 ? _GEN_2268 : _GEN_1244; // @[Sbuffer.scala 134:17]
  wire  _GEN_3293 = line_mask_clean_valid_1 ? _GEN_2269 : _GEN_1245; // @[Sbuffer.scala 134:17]
  wire  _GEN_3294 = line_mask_clean_valid_1 ? _GEN_2270 : _GEN_1246; // @[Sbuffer.scala 134:17]
  wire  _GEN_3295 = line_mask_clean_valid_1 ? _GEN_2271 : _GEN_1247; // @[Sbuffer.scala 134:17]
  wire  _GEN_3296 = line_mask_clean_valid_1 ? _GEN_2272 : _GEN_1248; // @[Sbuffer.scala 134:17]
  wire  _GEN_3297 = line_mask_clean_valid_1 ? _GEN_2273 : _GEN_1249; // @[Sbuffer.scala 134:17]
  wire  _GEN_3298 = line_mask_clean_valid_1 ? _GEN_2274 : _GEN_1250; // @[Sbuffer.scala 134:17]
  wire  _GEN_3299 = line_mask_clean_valid_1 ? _GEN_2275 : _GEN_1251; // @[Sbuffer.scala 134:17]
  wire  _GEN_3300 = line_mask_clean_valid_1 ? _GEN_2276 : _GEN_1252; // @[Sbuffer.scala 134:17]
  wire  _GEN_3301 = line_mask_clean_valid_1 ? _GEN_2277 : _GEN_1253; // @[Sbuffer.scala 134:17]
  wire  _GEN_3302 = line_mask_clean_valid_1 ? _GEN_2278 : _GEN_1254; // @[Sbuffer.scala 134:17]
  wire  _GEN_3303 = line_mask_clean_valid_1 ? _GEN_2279 : _GEN_1255; // @[Sbuffer.scala 134:17]
  wire  _GEN_3304 = line_mask_clean_valid_1 ? _GEN_2280 : _GEN_1256; // @[Sbuffer.scala 134:17]
  wire  _GEN_3305 = line_mask_clean_valid_1 ? _GEN_2281 : _GEN_1257; // @[Sbuffer.scala 134:17]
  wire  _GEN_3306 = line_mask_clean_valid_1 ? _GEN_2282 : _GEN_1258; // @[Sbuffer.scala 134:17]
  wire  _GEN_3307 = line_mask_clean_valid_1 ? _GEN_2283 : _GEN_1259; // @[Sbuffer.scala 134:17]
  wire  _GEN_3308 = line_mask_clean_valid_1 ? _GEN_2284 : _GEN_1260; // @[Sbuffer.scala 134:17]
  wire  _GEN_3309 = line_mask_clean_valid_1 ? _GEN_2285 : _GEN_1261; // @[Sbuffer.scala 134:17]
  wire  _GEN_3310 = line_mask_clean_valid_1 ? _GEN_2286 : _GEN_1262; // @[Sbuffer.scala 134:17]
  wire  _GEN_3311 = line_mask_clean_valid_1 ? _GEN_2287 : _GEN_1263; // @[Sbuffer.scala 134:17]
  wire  _GEN_3312 = line_mask_clean_valid_1 ? _GEN_2288 : _GEN_1264; // @[Sbuffer.scala 134:17]
  wire  _GEN_3313 = line_mask_clean_valid_1 ? _GEN_2289 : _GEN_1265; // @[Sbuffer.scala 134:17]
  wire  _GEN_3314 = line_mask_clean_valid_1 ? _GEN_2290 : _GEN_1266; // @[Sbuffer.scala 134:17]
  wire  _GEN_3315 = line_mask_clean_valid_1 ? _GEN_2291 : _GEN_1267; // @[Sbuffer.scala 134:17]
  wire  _GEN_3316 = line_mask_clean_valid_1 ? _GEN_2292 : _GEN_1268; // @[Sbuffer.scala 134:17]
  wire  _GEN_3317 = line_mask_clean_valid_1 ? _GEN_2293 : _GEN_1269; // @[Sbuffer.scala 134:17]
  wire  _GEN_3318 = line_mask_clean_valid_1 ? _GEN_2294 : _GEN_1270; // @[Sbuffer.scala 134:17]
  wire  _GEN_3319 = line_mask_clean_valid_1 ? _GEN_2295 : _GEN_1271; // @[Sbuffer.scala 134:17]
  wire  _GEN_3320 = line_mask_clean_valid_1 ? _GEN_2296 : _GEN_1272; // @[Sbuffer.scala 134:17]
  wire  _GEN_3321 = line_mask_clean_valid_1 ? _GEN_2297 : _GEN_1273; // @[Sbuffer.scala 134:17]
  wire  _GEN_3322 = line_mask_clean_valid_1 ? _GEN_2298 : _GEN_1274; // @[Sbuffer.scala 134:17]
  wire  _GEN_3323 = line_mask_clean_valid_1 ? _GEN_2299 : _GEN_1275; // @[Sbuffer.scala 134:17]
  wire  _GEN_3324 = line_mask_clean_valid_1 ? _GEN_2300 : _GEN_1276; // @[Sbuffer.scala 134:17]
  wire  _GEN_3325 = line_mask_clean_valid_1 ? _GEN_2301 : _GEN_1277; // @[Sbuffer.scala 134:17]
  wire  _GEN_3326 = line_mask_clean_valid_1 ? _GEN_2302 : _GEN_1278; // @[Sbuffer.scala 134:17]
  wire  _GEN_3327 = line_mask_clean_valid_1 ? _GEN_2303 : _GEN_1279; // @[Sbuffer.scala 134:17]
  wire  _GEN_3328 = line_mask_clean_valid_1 ? _GEN_2304 : _GEN_1280; // @[Sbuffer.scala 134:17]
  wire  _GEN_3329 = line_mask_clean_valid_1 ? _GEN_2305 : _GEN_1281; // @[Sbuffer.scala 134:17]
  wire  _GEN_3330 = line_mask_clean_valid_1 ? _GEN_2306 : _GEN_1282; // @[Sbuffer.scala 134:17]
  wire  _GEN_3331 = line_mask_clean_valid_1 ? _GEN_2307 : _GEN_1283; // @[Sbuffer.scala 134:17]
  wire  _GEN_3332 = line_mask_clean_valid_1 ? _GEN_2308 : _GEN_1284; // @[Sbuffer.scala 134:17]
  wire  _GEN_3333 = line_mask_clean_valid_1 ? _GEN_2309 : _GEN_1285; // @[Sbuffer.scala 134:17]
  wire  _GEN_3334 = line_mask_clean_valid_1 ? _GEN_2310 : _GEN_1286; // @[Sbuffer.scala 134:17]
  wire  _GEN_3335 = line_mask_clean_valid_1 ? _GEN_2311 : _GEN_1287; // @[Sbuffer.scala 134:17]
  wire  _GEN_3336 = line_mask_clean_valid_1 ? _GEN_2312 : _GEN_1288; // @[Sbuffer.scala 134:17]
  wire  _GEN_3337 = line_mask_clean_valid_1 ? _GEN_2313 : _GEN_1289; // @[Sbuffer.scala 134:17]
  wire  _GEN_3338 = line_mask_clean_valid_1 ? _GEN_2314 : _GEN_1290; // @[Sbuffer.scala 134:17]
  wire  _GEN_3339 = line_mask_clean_valid_1 ? _GEN_2315 : _GEN_1291; // @[Sbuffer.scala 134:17]
  wire  _GEN_3340 = line_mask_clean_valid_1 ? _GEN_2316 : _GEN_1292; // @[Sbuffer.scala 134:17]
  wire  _GEN_3341 = line_mask_clean_valid_1 ? _GEN_2317 : _GEN_1293; // @[Sbuffer.scala 134:17]
  wire  _GEN_3342 = line_mask_clean_valid_1 ? _GEN_2318 : _GEN_1294; // @[Sbuffer.scala 134:17]
  wire  _GEN_3343 = line_mask_clean_valid_1 ? _GEN_2319 : _GEN_1295; // @[Sbuffer.scala 134:17]
  wire  _GEN_3344 = line_mask_clean_valid_1 ? _GEN_2320 : _GEN_1296; // @[Sbuffer.scala 134:17]
  wire  _GEN_3345 = line_mask_clean_valid_1 ? _GEN_2321 : _GEN_1297; // @[Sbuffer.scala 134:17]
  wire  _GEN_3346 = line_mask_clean_valid_1 ? _GEN_2322 : _GEN_1298; // @[Sbuffer.scala 134:17]
  wire  _GEN_3347 = line_mask_clean_valid_1 ? _GEN_2323 : _GEN_1299; // @[Sbuffer.scala 134:17]
  wire  _GEN_3348 = line_mask_clean_valid_1 ? _GEN_2324 : _GEN_1300; // @[Sbuffer.scala 134:17]
  wire  _GEN_3349 = line_mask_clean_valid_1 ? _GEN_2325 : _GEN_1301; // @[Sbuffer.scala 134:17]
  wire  _GEN_3350 = line_mask_clean_valid_1 ? _GEN_2326 : _GEN_1302; // @[Sbuffer.scala 134:17]
  wire  _GEN_3351 = line_mask_clean_valid_1 ? _GEN_2327 : _GEN_1303; // @[Sbuffer.scala 134:17]
  wire  _GEN_3352 = line_mask_clean_valid_1 ? _GEN_2328 : _GEN_1304; // @[Sbuffer.scala 134:17]
  wire  _GEN_3353 = line_mask_clean_valid_1 ? _GEN_2329 : _GEN_1305; // @[Sbuffer.scala 134:17]
  wire  _GEN_3354 = line_mask_clean_valid_1 ? _GEN_2330 : _GEN_1306; // @[Sbuffer.scala 134:17]
  wire  _GEN_3355 = line_mask_clean_valid_1 ? _GEN_2331 : _GEN_1307; // @[Sbuffer.scala 134:17]
  wire  _GEN_3356 = line_mask_clean_valid_1 ? _GEN_2332 : _GEN_1308; // @[Sbuffer.scala 134:17]
  wire  _GEN_3357 = line_mask_clean_valid_1 ? _GEN_2333 : _GEN_1309; // @[Sbuffer.scala 134:17]
  wire  _GEN_3358 = line_mask_clean_valid_1 ? _GEN_2334 : _GEN_1310; // @[Sbuffer.scala 134:17]
  wire  _GEN_3359 = line_mask_clean_valid_1 ? _GEN_2335 : _GEN_1311; // @[Sbuffer.scala 134:17]
  wire  _GEN_3360 = line_mask_clean_valid_1 ? _GEN_2336 : _GEN_1312; // @[Sbuffer.scala 134:17]
  wire  _GEN_3361 = line_mask_clean_valid_1 ? _GEN_2337 : _GEN_1313; // @[Sbuffer.scala 134:17]
  wire  _GEN_3362 = line_mask_clean_valid_1 ? _GEN_2338 : _GEN_1314; // @[Sbuffer.scala 134:17]
  wire  _GEN_3363 = line_mask_clean_valid_1 ? _GEN_2339 : _GEN_1315; // @[Sbuffer.scala 134:17]
  wire  _GEN_3364 = line_mask_clean_valid_1 ? _GEN_2340 : _GEN_1316; // @[Sbuffer.scala 134:17]
  wire  _GEN_3365 = line_mask_clean_valid_1 ? _GEN_2341 : _GEN_1317; // @[Sbuffer.scala 134:17]
  wire  _GEN_3366 = line_mask_clean_valid_1 ? _GEN_2342 : _GEN_1318; // @[Sbuffer.scala 134:17]
  wire  _GEN_3367 = line_mask_clean_valid_1 ? _GEN_2343 : _GEN_1319; // @[Sbuffer.scala 134:17]
  wire  _GEN_3368 = line_mask_clean_valid_1 ? _GEN_2344 : _GEN_1320; // @[Sbuffer.scala 134:17]
  wire  _GEN_3369 = line_mask_clean_valid_1 ? _GEN_2345 : _GEN_1321; // @[Sbuffer.scala 134:17]
  wire  _GEN_3370 = line_mask_clean_valid_1 ? _GEN_2346 : _GEN_1322; // @[Sbuffer.scala 134:17]
  wire  _GEN_3371 = line_mask_clean_valid_1 ? _GEN_2347 : _GEN_1323; // @[Sbuffer.scala 134:17]
  wire  _GEN_3372 = line_mask_clean_valid_1 ? _GEN_2348 : _GEN_1324; // @[Sbuffer.scala 134:17]
  wire  _GEN_3373 = line_mask_clean_valid_1 ? _GEN_2349 : _GEN_1325; // @[Sbuffer.scala 134:17]
  wire  _GEN_3374 = line_mask_clean_valid_1 ? _GEN_2350 : _GEN_1326; // @[Sbuffer.scala 134:17]
  wire  _GEN_3375 = line_mask_clean_valid_1 ? _GEN_2351 : _GEN_1327; // @[Sbuffer.scala 134:17]
  wire  _GEN_3376 = line_mask_clean_valid_1 ? _GEN_2352 : _GEN_1328; // @[Sbuffer.scala 134:17]
  wire  _GEN_3377 = line_mask_clean_valid_1 ? _GEN_2353 : _GEN_1329; // @[Sbuffer.scala 134:17]
  wire  _GEN_3378 = line_mask_clean_valid_1 ? _GEN_2354 : _GEN_1330; // @[Sbuffer.scala 134:17]
  wire  _GEN_3379 = line_mask_clean_valid_1 ? _GEN_2355 : _GEN_1331; // @[Sbuffer.scala 134:17]
  wire  _GEN_3380 = line_mask_clean_valid_1 ? _GEN_2356 : _GEN_1332; // @[Sbuffer.scala 134:17]
  wire  _GEN_3381 = line_mask_clean_valid_1 ? _GEN_2357 : _GEN_1333; // @[Sbuffer.scala 134:17]
  wire  _GEN_3382 = line_mask_clean_valid_1 ? _GEN_2358 : _GEN_1334; // @[Sbuffer.scala 134:17]
  wire  _GEN_3383 = line_mask_clean_valid_1 ? _GEN_2359 : _GEN_1335; // @[Sbuffer.scala 134:17]
  wire  _GEN_3384 = line_mask_clean_valid_1 ? _GEN_2360 : _GEN_1336; // @[Sbuffer.scala 134:17]
  wire  _GEN_3385 = line_mask_clean_valid_1 ? _GEN_2361 : _GEN_1337; // @[Sbuffer.scala 134:17]
  wire  _GEN_3386 = line_mask_clean_valid_1 ? _GEN_2362 : _GEN_1338; // @[Sbuffer.scala 134:17]
  wire  _GEN_3387 = line_mask_clean_valid_1 ? _GEN_2363 : _GEN_1339; // @[Sbuffer.scala 134:17]
  wire  _GEN_3388 = line_mask_clean_valid_1 ? _GEN_2364 : _GEN_1340; // @[Sbuffer.scala 134:17]
  wire  _GEN_3389 = line_mask_clean_valid_1 ? _GEN_2365 : _GEN_1341; // @[Sbuffer.scala 134:17]
  wire  _GEN_3390 = line_mask_clean_valid_1 ? _GEN_2366 : _GEN_1342; // @[Sbuffer.scala 134:17]
  wire  _GEN_3391 = line_mask_clean_valid_1 ? _GEN_2367 : _GEN_1343; // @[Sbuffer.scala 134:17]
  wire  _GEN_3392 = line_mask_clean_valid_1 ? _GEN_2368 : _GEN_1344; // @[Sbuffer.scala 134:17]
  wire  _GEN_3393 = line_mask_clean_valid_1 ? _GEN_2369 : _GEN_1345; // @[Sbuffer.scala 134:17]
  wire  _GEN_3394 = line_mask_clean_valid_1 ? _GEN_2370 : _GEN_1346; // @[Sbuffer.scala 134:17]
  wire  _GEN_3395 = line_mask_clean_valid_1 ? _GEN_2371 : _GEN_1347; // @[Sbuffer.scala 134:17]
  wire  _GEN_3396 = line_mask_clean_valid_1 ? _GEN_2372 : _GEN_1348; // @[Sbuffer.scala 134:17]
  wire  _GEN_3397 = line_mask_clean_valid_1 ? _GEN_2373 : _GEN_1349; // @[Sbuffer.scala 134:17]
  wire  _GEN_3398 = line_mask_clean_valid_1 ? _GEN_2374 : _GEN_1350; // @[Sbuffer.scala 134:17]
  wire  _GEN_3399 = line_mask_clean_valid_1 ? _GEN_2375 : _GEN_1351; // @[Sbuffer.scala 134:17]
  wire  _GEN_3400 = line_mask_clean_valid_1 ? _GEN_2376 : _GEN_1352; // @[Sbuffer.scala 134:17]
  wire  _GEN_3401 = line_mask_clean_valid_1 ? _GEN_2377 : _GEN_1353; // @[Sbuffer.scala 134:17]
  wire  _GEN_3402 = line_mask_clean_valid_1 ? _GEN_2378 : _GEN_1354; // @[Sbuffer.scala 134:17]
  wire  _GEN_3403 = line_mask_clean_valid_1 ? _GEN_2379 : _GEN_1355; // @[Sbuffer.scala 134:17]
  wire  _GEN_3404 = line_mask_clean_valid_1 ? _GEN_2380 : _GEN_1356; // @[Sbuffer.scala 134:17]
  wire  _GEN_3405 = line_mask_clean_valid_1 ? _GEN_2381 : _GEN_1357; // @[Sbuffer.scala 134:17]
  wire  _GEN_3406 = line_mask_clean_valid_1 ? _GEN_2382 : _GEN_1358; // @[Sbuffer.scala 134:17]
  wire  _GEN_3407 = line_mask_clean_valid_1 ? _GEN_2383 : _GEN_1359; // @[Sbuffer.scala 134:17]
  wire  _GEN_3408 = line_mask_clean_valid_1 ? _GEN_2384 : _GEN_1360; // @[Sbuffer.scala 134:17]
  wire  _GEN_3409 = line_mask_clean_valid_1 ? _GEN_2385 : _GEN_1361; // @[Sbuffer.scala 134:17]
  wire  _GEN_3410 = line_mask_clean_valid_1 ? _GEN_2386 : _GEN_1362; // @[Sbuffer.scala 134:17]
  wire  _GEN_3411 = line_mask_clean_valid_1 ? _GEN_2387 : _GEN_1363; // @[Sbuffer.scala 134:17]
  wire  _GEN_3412 = line_mask_clean_valid_1 ? _GEN_2388 : _GEN_1364; // @[Sbuffer.scala 134:17]
  wire  _GEN_3413 = line_mask_clean_valid_1 ? _GEN_2389 : _GEN_1365; // @[Sbuffer.scala 134:17]
  wire  _GEN_3414 = line_mask_clean_valid_1 ? _GEN_2390 : _GEN_1366; // @[Sbuffer.scala 134:17]
  wire  _GEN_3415 = line_mask_clean_valid_1 ? _GEN_2391 : _GEN_1367; // @[Sbuffer.scala 134:17]
  wire  _GEN_3416 = line_mask_clean_valid_1 ? _GEN_2392 : _GEN_1368; // @[Sbuffer.scala 134:17]
  wire  _GEN_3417 = line_mask_clean_valid_1 ? _GEN_2393 : _GEN_1369; // @[Sbuffer.scala 134:17]
  wire  _GEN_3418 = line_mask_clean_valid_1 ? _GEN_2394 : _GEN_1370; // @[Sbuffer.scala 134:17]
  wire  _GEN_3419 = line_mask_clean_valid_1 ? _GEN_2395 : _GEN_1371; // @[Sbuffer.scala 134:17]
  wire  _GEN_3420 = line_mask_clean_valid_1 ? _GEN_2396 : _GEN_1372; // @[Sbuffer.scala 134:17]
  wire  _GEN_3421 = line_mask_clean_valid_1 ? _GEN_2397 : _GEN_1373; // @[Sbuffer.scala 134:17]
  wire  _GEN_3422 = line_mask_clean_valid_1 ? _GEN_2398 : _GEN_1374; // @[Sbuffer.scala 134:17]
  wire  _GEN_3423 = line_mask_clean_valid_1 ? _GEN_2399 : _GEN_1375; // @[Sbuffer.scala 134:17]
  wire  _GEN_3424 = line_mask_clean_valid_1 ? _GEN_2400 : _GEN_1376; // @[Sbuffer.scala 134:17]
  wire  _GEN_3425 = line_mask_clean_valid_1 ? _GEN_2401 : _GEN_1377; // @[Sbuffer.scala 134:17]
  wire  _GEN_3426 = line_mask_clean_valid_1 ? _GEN_2402 : _GEN_1378; // @[Sbuffer.scala 134:17]
  wire  _GEN_3427 = line_mask_clean_valid_1 ? _GEN_2403 : _GEN_1379; // @[Sbuffer.scala 134:17]
  wire  _GEN_3428 = line_mask_clean_valid_1 ? _GEN_2404 : _GEN_1380; // @[Sbuffer.scala 134:17]
  wire  _GEN_3429 = line_mask_clean_valid_1 ? _GEN_2405 : _GEN_1381; // @[Sbuffer.scala 134:17]
  wire  _GEN_3430 = line_mask_clean_valid_1 ? _GEN_2406 : _GEN_1382; // @[Sbuffer.scala 134:17]
  wire  _GEN_3431 = line_mask_clean_valid_1 ? _GEN_2407 : _GEN_1383; // @[Sbuffer.scala 134:17]
  wire  _GEN_3432 = line_mask_clean_valid_1 ? _GEN_2408 : _GEN_1384; // @[Sbuffer.scala 134:17]
  wire  _GEN_3433 = line_mask_clean_valid_1 ? _GEN_2409 : _GEN_1385; // @[Sbuffer.scala 134:17]
  wire  _GEN_3434 = line_mask_clean_valid_1 ? _GEN_2410 : _GEN_1386; // @[Sbuffer.scala 134:17]
  wire  _GEN_3435 = line_mask_clean_valid_1 ? _GEN_2411 : _GEN_1387; // @[Sbuffer.scala 134:17]
  wire  _GEN_3436 = line_mask_clean_valid_1 ? _GEN_2412 : _GEN_1388; // @[Sbuffer.scala 134:17]
  wire  _GEN_3437 = line_mask_clean_valid_1 ? _GEN_2413 : _GEN_1389; // @[Sbuffer.scala 134:17]
  wire  _GEN_3438 = line_mask_clean_valid_1 ? _GEN_2414 : _GEN_1390; // @[Sbuffer.scala 134:17]
  wire  _GEN_3439 = line_mask_clean_valid_1 ? _GEN_2415 : _GEN_1391; // @[Sbuffer.scala 134:17]
  wire  _GEN_3440 = line_mask_clean_valid_1 ? _GEN_2416 : _GEN_1392; // @[Sbuffer.scala 134:17]
  wire  _GEN_3441 = line_mask_clean_valid_1 ? _GEN_2417 : _GEN_1393; // @[Sbuffer.scala 134:17]
  wire  _GEN_3442 = line_mask_clean_valid_1 ? _GEN_2418 : _GEN_1394; // @[Sbuffer.scala 134:17]
  wire  _GEN_3443 = line_mask_clean_valid_1 ? _GEN_2419 : _GEN_1395; // @[Sbuffer.scala 134:17]
  wire  _GEN_3444 = line_mask_clean_valid_1 ? _GEN_2420 : _GEN_1396; // @[Sbuffer.scala 134:17]
  wire  _GEN_3445 = line_mask_clean_valid_1 ? _GEN_2421 : _GEN_1397; // @[Sbuffer.scala 134:17]
  wire  _GEN_3446 = line_mask_clean_valid_1 ? _GEN_2422 : _GEN_1398; // @[Sbuffer.scala 134:17]
  wire  _GEN_3447 = line_mask_clean_valid_1 ? _GEN_2423 : _GEN_1399; // @[Sbuffer.scala 134:17]
  wire  _GEN_3448 = line_mask_clean_valid_1 ? _GEN_2424 : _GEN_1400; // @[Sbuffer.scala 134:17]
  wire  _GEN_3449 = line_mask_clean_valid_1 ? _GEN_2425 : _GEN_1401; // @[Sbuffer.scala 134:17]
  wire  _GEN_3450 = line_mask_clean_valid_1 ? _GEN_2426 : _GEN_1402; // @[Sbuffer.scala 134:17]
  wire  _GEN_3451 = line_mask_clean_valid_1 ? _GEN_2427 : _GEN_1403; // @[Sbuffer.scala 134:17]
  wire  _GEN_3452 = line_mask_clean_valid_1 ? _GEN_2428 : _GEN_1404; // @[Sbuffer.scala 134:17]
  wire  _GEN_3453 = line_mask_clean_valid_1 ? _GEN_2429 : _GEN_1405; // @[Sbuffer.scala 134:17]
  wire  _GEN_3454 = line_mask_clean_valid_1 ? _GEN_2430 : _GEN_1406; // @[Sbuffer.scala 134:17]
  wire  _GEN_3455 = line_mask_clean_valid_1 ? _GEN_2431 : _GEN_1407; // @[Sbuffer.scala 134:17]
  wire  _GEN_3456 = line_mask_clean_valid_1 ? _GEN_2432 : _GEN_1408; // @[Sbuffer.scala 134:17]
  wire  _GEN_3457 = line_mask_clean_valid_1 ? _GEN_2433 : _GEN_1409; // @[Sbuffer.scala 134:17]
  wire  _GEN_3458 = line_mask_clean_valid_1 ? _GEN_2434 : _GEN_1410; // @[Sbuffer.scala 134:17]
  wire  _GEN_3459 = line_mask_clean_valid_1 ? _GEN_2435 : _GEN_1411; // @[Sbuffer.scala 134:17]
  wire  _GEN_3460 = line_mask_clean_valid_1 ? _GEN_2436 : _GEN_1412; // @[Sbuffer.scala 134:17]
  wire  _GEN_3461 = line_mask_clean_valid_1 ? _GEN_2437 : _GEN_1413; // @[Sbuffer.scala 134:17]
  wire  _GEN_3462 = line_mask_clean_valid_1 ? _GEN_2438 : _GEN_1414; // @[Sbuffer.scala 134:17]
  wire  _GEN_3463 = line_mask_clean_valid_1 ? _GEN_2439 : _GEN_1415; // @[Sbuffer.scala 134:17]
  wire  _GEN_3464 = line_mask_clean_valid_1 ? _GEN_2440 : _GEN_1416; // @[Sbuffer.scala 134:17]
  wire  _GEN_3465 = line_mask_clean_valid_1 ? _GEN_2441 : _GEN_1417; // @[Sbuffer.scala 134:17]
  wire  _GEN_3466 = line_mask_clean_valid_1 ? _GEN_2442 : _GEN_1418; // @[Sbuffer.scala 134:17]
  wire  _GEN_3467 = line_mask_clean_valid_1 ? _GEN_2443 : _GEN_1419; // @[Sbuffer.scala 134:17]
  wire  _GEN_3468 = line_mask_clean_valid_1 ? _GEN_2444 : _GEN_1420; // @[Sbuffer.scala 134:17]
  wire  _GEN_3469 = line_mask_clean_valid_1 ? _GEN_2445 : _GEN_1421; // @[Sbuffer.scala 134:17]
  wire  _GEN_3470 = line_mask_clean_valid_1 ? _GEN_2446 : _GEN_1422; // @[Sbuffer.scala 134:17]
  wire  _GEN_3471 = line_mask_clean_valid_1 ? _GEN_2447 : _GEN_1423; // @[Sbuffer.scala 134:17]
  wire  _GEN_3472 = line_mask_clean_valid_1 ? _GEN_2448 : _GEN_1424; // @[Sbuffer.scala 134:17]
  wire  _GEN_3473 = line_mask_clean_valid_1 ? _GEN_2449 : _GEN_1425; // @[Sbuffer.scala 134:17]
  wire  _GEN_3474 = line_mask_clean_valid_1 ? _GEN_2450 : _GEN_1426; // @[Sbuffer.scala 134:17]
  wire  _GEN_3475 = line_mask_clean_valid_1 ? _GEN_2451 : _GEN_1427; // @[Sbuffer.scala 134:17]
  wire  _GEN_3476 = line_mask_clean_valid_1 ? _GEN_2452 : _GEN_1428; // @[Sbuffer.scala 134:17]
  wire  _GEN_3477 = line_mask_clean_valid_1 ? _GEN_2453 : _GEN_1429; // @[Sbuffer.scala 134:17]
  wire  _GEN_3478 = line_mask_clean_valid_1 ? _GEN_2454 : _GEN_1430; // @[Sbuffer.scala 134:17]
  wire  _GEN_3479 = line_mask_clean_valid_1 ? _GEN_2455 : _GEN_1431; // @[Sbuffer.scala 134:17]
  wire  _GEN_3480 = line_mask_clean_valid_1 ? _GEN_2456 : _GEN_1432; // @[Sbuffer.scala 134:17]
  wire  _GEN_3481 = line_mask_clean_valid_1 ? _GEN_2457 : _GEN_1433; // @[Sbuffer.scala 134:17]
  wire  _GEN_3482 = line_mask_clean_valid_1 ? _GEN_2458 : _GEN_1434; // @[Sbuffer.scala 134:17]
  wire  _GEN_3483 = line_mask_clean_valid_1 ? _GEN_2459 : _GEN_1435; // @[Sbuffer.scala 134:17]
  wire  _GEN_3484 = line_mask_clean_valid_1 ? _GEN_2460 : _GEN_1436; // @[Sbuffer.scala 134:17]
  wire  _GEN_3485 = line_mask_clean_valid_1 ? _GEN_2461 : _GEN_1437; // @[Sbuffer.scala 134:17]
  wire  _GEN_3486 = line_mask_clean_valid_1 ? _GEN_2462 : _GEN_1438; // @[Sbuffer.scala 134:17]
  wire  _GEN_3487 = line_mask_clean_valid_1 ? _GEN_2463 : _GEN_1439; // @[Sbuffer.scala 134:17]
  wire  _GEN_3488 = line_mask_clean_valid_1 ? _GEN_2464 : _GEN_1440; // @[Sbuffer.scala 134:17]
  wire  _GEN_3489 = line_mask_clean_valid_1 ? _GEN_2465 : _GEN_1441; // @[Sbuffer.scala 134:17]
  wire  _GEN_3490 = line_mask_clean_valid_1 ? _GEN_2466 : _GEN_1442; // @[Sbuffer.scala 134:17]
  wire  _GEN_3491 = line_mask_clean_valid_1 ? _GEN_2467 : _GEN_1443; // @[Sbuffer.scala 134:17]
  wire  _GEN_3492 = line_mask_clean_valid_1 ? _GEN_2468 : _GEN_1444; // @[Sbuffer.scala 134:17]
  wire  _GEN_3493 = line_mask_clean_valid_1 ? _GEN_2469 : _GEN_1445; // @[Sbuffer.scala 134:17]
  wire  _GEN_3494 = line_mask_clean_valid_1 ? _GEN_2470 : _GEN_1446; // @[Sbuffer.scala 134:17]
  wire  _GEN_3495 = line_mask_clean_valid_1 ? _GEN_2471 : _GEN_1447; // @[Sbuffer.scala 134:17]
  wire  _GEN_3496 = line_mask_clean_valid_1 ? _GEN_2472 : _GEN_1448; // @[Sbuffer.scala 134:17]
  wire  _GEN_3497 = line_mask_clean_valid_1 ? _GEN_2473 : _GEN_1449; // @[Sbuffer.scala 134:17]
  wire  _GEN_3498 = line_mask_clean_valid_1 ? _GEN_2474 : _GEN_1450; // @[Sbuffer.scala 134:17]
  wire  _GEN_3499 = line_mask_clean_valid_1 ? _GEN_2475 : _GEN_1451; // @[Sbuffer.scala 134:17]
  wire  _GEN_3500 = line_mask_clean_valid_1 ? _GEN_2476 : _GEN_1452; // @[Sbuffer.scala 134:17]
  wire  _GEN_3501 = line_mask_clean_valid_1 ? _GEN_2477 : _GEN_1453; // @[Sbuffer.scala 134:17]
  wire  _GEN_3502 = line_mask_clean_valid_1 ? _GEN_2478 : _GEN_1454; // @[Sbuffer.scala 134:17]
  wire  _GEN_3503 = line_mask_clean_valid_1 ? _GEN_2479 : _GEN_1455; // @[Sbuffer.scala 134:17]
  wire  _GEN_3504 = line_mask_clean_valid_1 ? _GEN_2480 : _GEN_1456; // @[Sbuffer.scala 134:17]
  wire  _GEN_3505 = line_mask_clean_valid_1 ? _GEN_2481 : _GEN_1457; // @[Sbuffer.scala 134:17]
  wire  _GEN_3506 = line_mask_clean_valid_1 ? _GEN_2482 : _GEN_1458; // @[Sbuffer.scala 134:17]
  wire  _GEN_3507 = line_mask_clean_valid_1 ? _GEN_2483 : _GEN_1459; // @[Sbuffer.scala 134:17]
  wire  _GEN_3508 = line_mask_clean_valid_1 ? _GEN_2484 : _GEN_1460; // @[Sbuffer.scala 134:17]
  wire  _GEN_3509 = line_mask_clean_valid_1 ? _GEN_2485 : _GEN_1461; // @[Sbuffer.scala 134:17]
  wire  _GEN_3510 = line_mask_clean_valid_1 ? _GEN_2486 : _GEN_1462; // @[Sbuffer.scala 134:17]
  wire  _GEN_3511 = line_mask_clean_valid_1 ? _GEN_2487 : _GEN_1463; // @[Sbuffer.scala 134:17]
  wire  _GEN_3512 = line_mask_clean_valid_1 ? _GEN_2488 : _GEN_1464; // @[Sbuffer.scala 134:17]
  wire  _GEN_3513 = line_mask_clean_valid_1 ? _GEN_2489 : _GEN_1465; // @[Sbuffer.scala 134:17]
  wire  _GEN_3514 = line_mask_clean_valid_1 ? _GEN_2490 : _GEN_1466; // @[Sbuffer.scala 134:17]
  wire  _GEN_3515 = line_mask_clean_valid_1 ? _GEN_2491 : _GEN_1467; // @[Sbuffer.scala 134:17]
  wire  _GEN_3516 = line_mask_clean_valid_1 ? _GEN_2492 : _GEN_1468; // @[Sbuffer.scala 134:17]
  wire  _GEN_3517 = line_mask_clean_valid_1 ? _GEN_2493 : _GEN_1469; // @[Sbuffer.scala 134:17]
  wire  _GEN_3518 = line_mask_clean_valid_1 ? _GEN_2494 : _GEN_1470; // @[Sbuffer.scala 134:17]
  wire  _GEN_3519 = line_mask_clean_valid_1 ? _GEN_2495 : _GEN_1471; // @[Sbuffer.scala 134:17]
  wire  _GEN_3520 = line_mask_clean_valid_1 ? _GEN_2496 : _GEN_1472; // @[Sbuffer.scala 134:17]
  wire  _GEN_3521 = line_mask_clean_valid_1 ? _GEN_2497 : _GEN_1473; // @[Sbuffer.scala 134:17]
  wire  _GEN_3522 = line_mask_clean_valid_1 ? _GEN_2498 : _GEN_1474; // @[Sbuffer.scala 134:17]
  wire  _GEN_3523 = line_mask_clean_valid_1 ? _GEN_2499 : _GEN_1475; // @[Sbuffer.scala 134:17]
  wire  _GEN_3524 = line_mask_clean_valid_1 ? _GEN_2500 : _GEN_1476; // @[Sbuffer.scala 134:17]
  wire  _GEN_3525 = line_mask_clean_valid_1 ? _GEN_2501 : _GEN_1477; // @[Sbuffer.scala 134:17]
  wire  _GEN_3526 = line_mask_clean_valid_1 ? _GEN_2502 : _GEN_1478; // @[Sbuffer.scala 134:17]
  wire  _GEN_3527 = line_mask_clean_valid_1 ? _GEN_2503 : _GEN_1479; // @[Sbuffer.scala 134:17]
  wire  _GEN_3528 = line_mask_clean_valid_1 ? _GEN_2504 : _GEN_1480; // @[Sbuffer.scala 134:17]
  wire  _GEN_3529 = line_mask_clean_valid_1 ? _GEN_2505 : _GEN_1481; // @[Sbuffer.scala 134:17]
  wire  _GEN_3530 = line_mask_clean_valid_1 ? _GEN_2506 : _GEN_1482; // @[Sbuffer.scala 134:17]
  wire  _GEN_3531 = line_mask_clean_valid_1 ? _GEN_2507 : _GEN_1483; // @[Sbuffer.scala 134:17]
  wire  _GEN_3532 = line_mask_clean_valid_1 ? _GEN_2508 : _GEN_1484; // @[Sbuffer.scala 134:17]
  wire  _GEN_3533 = line_mask_clean_valid_1 ? _GEN_2509 : _GEN_1485; // @[Sbuffer.scala 134:17]
  wire  _GEN_3534 = line_mask_clean_valid_1 ? _GEN_2510 : _GEN_1486; // @[Sbuffer.scala 134:17]
  wire  _GEN_3535 = line_mask_clean_valid_1 ? _GEN_2511 : _GEN_1487; // @[Sbuffer.scala 134:17]
  wire  _GEN_3536 = line_mask_clean_valid_1 ? _GEN_2512 : _GEN_1488; // @[Sbuffer.scala 134:17]
  wire  _GEN_3537 = line_mask_clean_valid_1 ? _GEN_2513 : _GEN_1489; // @[Sbuffer.scala 134:17]
  wire  _GEN_3538 = line_mask_clean_valid_1 ? _GEN_2514 : _GEN_1490; // @[Sbuffer.scala 134:17]
  wire  _GEN_3539 = line_mask_clean_valid_1 ? _GEN_2515 : _GEN_1491; // @[Sbuffer.scala 134:17]
  wire  _GEN_3540 = line_mask_clean_valid_1 ? _GEN_2516 : _GEN_1492; // @[Sbuffer.scala 134:17]
  wire  _GEN_3541 = line_mask_clean_valid_1 ? _GEN_2517 : _GEN_1493; // @[Sbuffer.scala 134:17]
  wire  _GEN_3542 = line_mask_clean_valid_1 ? _GEN_2518 : _GEN_1494; // @[Sbuffer.scala 134:17]
  wire  _GEN_3543 = line_mask_clean_valid_1 ? _GEN_2519 : _GEN_1495; // @[Sbuffer.scala 134:17]
  wire  _GEN_3544 = line_mask_clean_valid_1 ? _GEN_2520 : _GEN_1496; // @[Sbuffer.scala 134:17]
  wire  _GEN_3545 = line_mask_clean_valid_1 ? _GEN_2521 : _GEN_1497; // @[Sbuffer.scala 134:17]
  wire  _GEN_3546 = line_mask_clean_valid_1 ? _GEN_2522 : _GEN_1498; // @[Sbuffer.scala 134:17]
  wire  _GEN_3547 = line_mask_clean_valid_1 ? _GEN_2523 : _GEN_1499; // @[Sbuffer.scala 134:17]
  wire  _GEN_3548 = line_mask_clean_valid_1 ? _GEN_2524 : _GEN_1500; // @[Sbuffer.scala 134:17]
  wire  _GEN_3549 = line_mask_clean_valid_1 ? _GEN_2525 : _GEN_1501; // @[Sbuffer.scala 134:17]
  wire  _GEN_3550 = line_mask_clean_valid_1 ? _GEN_2526 : _GEN_1502; // @[Sbuffer.scala 134:17]
  wire  _GEN_3551 = line_mask_clean_valid_1 ? _GEN_2527 : _GEN_1503; // @[Sbuffer.scala 134:17]
  wire  _GEN_3552 = line_mask_clean_valid_1 ? _GEN_2528 : _GEN_1504; // @[Sbuffer.scala 134:17]
  wire  _GEN_3553 = line_mask_clean_valid_1 ? _GEN_2529 : _GEN_1505; // @[Sbuffer.scala 134:17]
  wire  _GEN_3554 = line_mask_clean_valid_1 ? _GEN_2530 : _GEN_1506; // @[Sbuffer.scala 134:17]
  wire  _GEN_3555 = line_mask_clean_valid_1 ? _GEN_2531 : _GEN_1507; // @[Sbuffer.scala 134:17]
  wire  _GEN_3556 = line_mask_clean_valid_1 ? _GEN_2532 : _GEN_1508; // @[Sbuffer.scala 134:17]
  wire  _GEN_3557 = line_mask_clean_valid_1 ? _GEN_2533 : _GEN_1509; // @[Sbuffer.scala 134:17]
  wire  _GEN_3558 = line_mask_clean_valid_1 ? _GEN_2534 : _GEN_1510; // @[Sbuffer.scala 134:17]
  wire  _GEN_3559 = line_mask_clean_valid_1 ? _GEN_2535 : _GEN_1511; // @[Sbuffer.scala 134:17]
  wire  _GEN_3560 = line_mask_clean_valid_1 ? _GEN_2536 : _GEN_1512; // @[Sbuffer.scala 134:17]
  wire  _GEN_3561 = line_mask_clean_valid_1 ? _GEN_2537 : _GEN_1513; // @[Sbuffer.scala 134:17]
  wire  _GEN_3562 = line_mask_clean_valid_1 ? _GEN_2538 : _GEN_1514; // @[Sbuffer.scala 134:17]
  wire  _GEN_3563 = line_mask_clean_valid_1 ? _GEN_2539 : _GEN_1515; // @[Sbuffer.scala 134:17]
  wire  _GEN_3564 = line_mask_clean_valid_1 ? _GEN_2540 : _GEN_1516; // @[Sbuffer.scala 134:17]
  wire  _GEN_3565 = line_mask_clean_valid_1 ? _GEN_2541 : _GEN_1517; // @[Sbuffer.scala 134:17]
  wire  _GEN_3566 = line_mask_clean_valid_1 ? _GEN_2542 : _GEN_1518; // @[Sbuffer.scala 134:17]
  wire  _GEN_3567 = line_mask_clean_valid_1 ? _GEN_2543 : _GEN_1519; // @[Sbuffer.scala 134:17]
  wire  _GEN_3568 = line_mask_clean_valid_1 ? _GEN_2544 : _GEN_1520; // @[Sbuffer.scala 134:17]
  wire  _GEN_3569 = line_mask_clean_valid_1 ? _GEN_2545 : _GEN_1521; // @[Sbuffer.scala 134:17]
  wire  _GEN_3570 = line_mask_clean_valid_1 ? _GEN_2546 : _GEN_1522; // @[Sbuffer.scala 134:17]
  wire  _GEN_3571 = line_mask_clean_valid_1 ? _GEN_2547 : _GEN_1523; // @[Sbuffer.scala 134:17]
  wire  _GEN_3572 = line_mask_clean_valid_1 ? _GEN_2548 : _GEN_1524; // @[Sbuffer.scala 134:17]
  wire  _GEN_3573 = line_mask_clean_valid_1 ? _GEN_2549 : _GEN_1525; // @[Sbuffer.scala 134:17]
  wire  _GEN_3574 = line_mask_clean_valid_1 ? _GEN_2550 : _GEN_1526; // @[Sbuffer.scala 134:17]
  wire  _GEN_3575 = line_mask_clean_valid_1 ? _GEN_2551 : _GEN_1527; // @[Sbuffer.scala 134:17]
  wire  _GEN_3576 = line_mask_clean_valid_1 ? _GEN_2552 : _GEN_1528; // @[Sbuffer.scala 134:17]
  wire  _GEN_3577 = line_mask_clean_valid_1 ? _GEN_2553 : _GEN_1529; // @[Sbuffer.scala 134:17]
  wire  _GEN_3578 = line_mask_clean_valid_1 ? _GEN_2554 : _GEN_1530; // @[Sbuffer.scala 134:17]
  wire  _GEN_3579 = line_mask_clean_valid_1 ? _GEN_2555 : _GEN_1531; // @[Sbuffer.scala 134:17]
  wire  _GEN_3580 = line_mask_clean_valid_1 ? _GEN_2556 : _GEN_1532; // @[Sbuffer.scala 134:17]
  wire  _GEN_3581 = line_mask_clean_valid_1 ? _GEN_2557 : _GEN_1533; // @[Sbuffer.scala 134:17]
  wire  _GEN_3582 = line_mask_clean_valid_1 ? _GEN_2558 : _GEN_1534; // @[Sbuffer.scala 134:17]
  wire  _GEN_3583 = line_mask_clean_valid_1 ? _GEN_2559 : _GEN_1535; // @[Sbuffer.scala 134:17]
  wire  _GEN_3584 = line_mask_clean_valid_1 ? _GEN_2560 : _GEN_1536; // @[Sbuffer.scala 134:17]
  wire  _GEN_3585 = line_mask_clean_valid_1 ? _GEN_2561 : _GEN_1537; // @[Sbuffer.scala 134:17]
  wire  _GEN_3586 = line_mask_clean_valid_1 ? _GEN_2562 : _GEN_1538; // @[Sbuffer.scala 134:17]
  wire  _GEN_3587 = line_mask_clean_valid_1 ? _GEN_2563 : _GEN_1539; // @[Sbuffer.scala 134:17]
  wire  _GEN_3588 = line_mask_clean_valid_1 ? _GEN_2564 : _GEN_1540; // @[Sbuffer.scala 134:17]
  wire  _GEN_3589 = line_mask_clean_valid_1 ? _GEN_2565 : _GEN_1541; // @[Sbuffer.scala 134:17]
  wire  _GEN_3590 = line_mask_clean_valid_1 ? _GEN_2566 : _GEN_1542; // @[Sbuffer.scala 134:17]
  wire  _GEN_3591 = line_mask_clean_valid_1 ? _GEN_2567 : _GEN_1543; // @[Sbuffer.scala 134:17]
  wire  _GEN_3592 = line_mask_clean_valid_1 ? _GEN_2568 : _GEN_1544; // @[Sbuffer.scala 134:17]
  wire  _GEN_3593 = line_mask_clean_valid_1 ? _GEN_2569 : _GEN_1545; // @[Sbuffer.scala 134:17]
  wire  _GEN_3594 = line_mask_clean_valid_1 ? _GEN_2570 : _GEN_1546; // @[Sbuffer.scala 134:17]
  wire  _GEN_3595 = line_mask_clean_valid_1 ? _GEN_2571 : _GEN_1547; // @[Sbuffer.scala 134:17]
  wire  _GEN_3596 = line_mask_clean_valid_1 ? _GEN_2572 : _GEN_1548; // @[Sbuffer.scala 134:17]
  wire  _GEN_3597 = line_mask_clean_valid_1 ? _GEN_2573 : _GEN_1549; // @[Sbuffer.scala 134:17]
  wire  _GEN_3598 = line_mask_clean_valid_1 ? _GEN_2574 : _GEN_1550; // @[Sbuffer.scala 134:17]
  wire  _GEN_3599 = line_mask_clean_valid_1 ? _GEN_2575 : _GEN_1551; // @[Sbuffer.scala 134:17]
  wire  _GEN_3600 = line_mask_clean_valid_1 ? _GEN_2576 : _GEN_1552; // @[Sbuffer.scala 134:17]
  wire  _GEN_3601 = line_mask_clean_valid_1 ? _GEN_2577 : _GEN_1553; // @[Sbuffer.scala 134:17]
  wire  _GEN_3602 = line_mask_clean_valid_1 ? _GEN_2578 : _GEN_1554; // @[Sbuffer.scala 134:17]
  wire  _GEN_3603 = line_mask_clean_valid_1 ? _GEN_2579 : _GEN_1555; // @[Sbuffer.scala 134:17]
  wire  _GEN_3604 = line_mask_clean_valid_1 ? _GEN_2580 : _GEN_1556; // @[Sbuffer.scala 134:17]
  wire  _GEN_3605 = line_mask_clean_valid_1 ? _GEN_2581 : _GEN_1557; // @[Sbuffer.scala 134:17]
  wire  _GEN_3606 = line_mask_clean_valid_1 ? _GEN_2582 : _GEN_1558; // @[Sbuffer.scala 134:17]
  wire  _GEN_3607 = line_mask_clean_valid_1 ? _GEN_2583 : _GEN_1559; // @[Sbuffer.scala 134:17]
  wire  _GEN_3608 = line_mask_clean_valid_1 ? _GEN_2584 : _GEN_1560; // @[Sbuffer.scala 134:17]
  wire  _GEN_3609 = line_mask_clean_valid_1 ? _GEN_2585 : _GEN_1561; // @[Sbuffer.scala 134:17]
  wire  _GEN_3610 = line_mask_clean_valid_1 ? _GEN_2586 : _GEN_1562; // @[Sbuffer.scala 134:17]
  wire  _GEN_3611 = line_mask_clean_valid_1 ? _GEN_2587 : _GEN_1563; // @[Sbuffer.scala 134:17]
  wire  _GEN_3612 = line_mask_clean_valid_1 ? _GEN_2588 : _GEN_1564; // @[Sbuffer.scala 134:17]
  wire  _GEN_3613 = line_mask_clean_valid_1 ? _GEN_2589 : _GEN_1565; // @[Sbuffer.scala 134:17]
  wire  _GEN_3614 = line_mask_clean_valid_1 ? _GEN_2590 : _GEN_1566; // @[Sbuffer.scala 134:17]
  wire  _GEN_3615 = line_mask_clean_valid_1 ? _GEN_2591 : _GEN_1567; // @[Sbuffer.scala 134:17]
  wire  _GEN_3616 = line_mask_clean_valid_1 ? _GEN_2592 : _GEN_1568; // @[Sbuffer.scala 134:17]
  wire  _GEN_3617 = line_mask_clean_valid_1 ? _GEN_2593 : _GEN_1569; // @[Sbuffer.scala 134:17]
  wire  _GEN_3618 = line_mask_clean_valid_1 ? _GEN_2594 : _GEN_1570; // @[Sbuffer.scala 134:17]
  wire  _GEN_3619 = line_mask_clean_valid_1 ? _GEN_2595 : _GEN_1571; // @[Sbuffer.scala 134:17]
  wire  _GEN_3620 = line_mask_clean_valid_1 ? _GEN_2596 : _GEN_1572; // @[Sbuffer.scala 134:17]
  wire  _GEN_3621 = line_mask_clean_valid_1 ? _GEN_2597 : _GEN_1573; // @[Sbuffer.scala 134:17]
  wire  _GEN_3622 = line_mask_clean_valid_1 ? _GEN_2598 : _GEN_1574; // @[Sbuffer.scala 134:17]
  wire  _GEN_3623 = line_mask_clean_valid_1 ? _GEN_2599 : _GEN_1575; // @[Sbuffer.scala 134:17]
  wire  _GEN_3624 = line_mask_clean_valid_1 ? _GEN_2600 : _GEN_1576; // @[Sbuffer.scala 134:17]
  wire  _GEN_3625 = line_mask_clean_valid_1 ? _GEN_2601 : _GEN_1577; // @[Sbuffer.scala 134:17]
  wire  _GEN_3626 = line_mask_clean_valid_1 ? _GEN_2602 : _GEN_1578; // @[Sbuffer.scala 134:17]
  wire  _GEN_3627 = line_mask_clean_valid_1 ? _GEN_2603 : _GEN_1579; // @[Sbuffer.scala 134:17]
  wire  _GEN_3628 = line_mask_clean_valid_1 ? _GEN_2604 : _GEN_1580; // @[Sbuffer.scala 134:17]
  wire  _GEN_3629 = line_mask_clean_valid_1 ? _GEN_2605 : _GEN_1581; // @[Sbuffer.scala 134:17]
  wire  _GEN_3630 = line_mask_clean_valid_1 ? _GEN_2606 : _GEN_1582; // @[Sbuffer.scala 134:17]
  wire  _GEN_3631 = line_mask_clean_valid_1 ? _GEN_2607 : _GEN_1583; // @[Sbuffer.scala 134:17]
  wire  _GEN_3632 = line_mask_clean_valid_1 ? _GEN_2608 : _GEN_1584; // @[Sbuffer.scala 134:17]
  wire  _GEN_3633 = line_mask_clean_valid_1 ? _GEN_2609 : _GEN_1585; // @[Sbuffer.scala 134:17]
  wire  _GEN_3634 = line_mask_clean_valid_1 ? _GEN_2610 : _GEN_1586; // @[Sbuffer.scala 134:17]
  wire  _GEN_3635 = line_mask_clean_valid_1 ? _GEN_2611 : _GEN_1587; // @[Sbuffer.scala 134:17]
  wire  _GEN_3636 = line_mask_clean_valid_1 ? _GEN_2612 : _GEN_1588; // @[Sbuffer.scala 134:17]
  wire  _GEN_3637 = line_mask_clean_valid_1 ? _GEN_2613 : _GEN_1589; // @[Sbuffer.scala 134:17]
  wire  _GEN_3638 = line_mask_clean_valid_1 ? _GEN_2614 : _GEN_1590; // @[Sbuffer.scala 134:17]
  wire  _GEN_3639 = line_mask_clean_valid_1 ? _GEN_2615 : _GEN_1591; // @[Sbuffer.scala 134:17]
  wire  _GEN_3640 = line_mask_clean_valid_1 ? _GEN_2616 : _GEN_1592; // @[Sbuffer.scala 134:17]
  wire  _GEN_3641 = line_mask_clean_valid_1 ? _GEN_2617 : _GEN_1593; // @[Sbuffer.scala 134:17]
  wire  _GEN_3642 = line_mask_clean_valid_1 ? _GEN_2618 : _GEN_1594; // @[Sbuffer.scala 134:17]
  wire  _GEN_3643 = line_mask_clean_valid_1 ? _GEN_2619 : _GEN_1595; // @[Sbuffer.scala 134:17]
  wire  _GEN_3644 = line_mask_clean_valid_1 ? _GEN_2620 : _GEN_1596; // @[Sbuffer.scala 134:17]
  wire  _GEN_3645 = line_mask_clean_valid_1 ? _GEN_2621 : _GEN_1597; // @[Sbuffer.scala 134:17]
  wire  _GEN_3646 = line_mask_clean_valid_1 ? _GEN_2622 : _GEN_1598; // @[Sbuffer.scala 134:17]
  wire  _GEN_3647 = line_mask_clean_valid_1 ? _GEN_2623 : _GEN_1599; // @[Sbuffer.scala 134:17]
  wire  _GEN_3648 = line_mask_clean_valid_1 ? _GEN_2624 : _GEN_1600; // @[Sbuffer.scala 134:17]
  wire  _GEN_3649 = line_mask_clean_valid_1 ? _GEN_2625 : _GEN_1601; // @[Sbuffer.scala 134:17]
  wire  _GEN_3650 = line_mask_clean_valid_1 ? _GEN_2626 : _GEN_1602; // @[Sbuffer.scala 134:17]
  wire  _GEN_3651 = line_mask_clean_valid_1 ? _GEN_2627 : _GEN_1603; // @[Sbuffer.scala 134:17]
  wire  _GEN_3652 = line_mask_clean_valid_1 ? _GEN_2628 : _GEN_1604; // @[Sbuffer.scala 134:17]
  wire  _GEN_3653 = line_mask_clean_valid_1 ? _GEN_2629 : _GEN_1605; // @[Sbuffer.scala 134:17]
  wire  _GEN_3654 = line_mask_clean_valid_1 ? _GEN_2630 : _GEN_1606; // @[Sbuffer.scala 134:17]
  wire  _GEN_3655 = line_mask_clean_valid_1 ? _GEN_2631 : _GEN_1607; // @[Sbuffer.scala 134:17]
  wire  _GEN_3656 = line_mask_clean_valid_1 ? _GEN_2632 : _GEN_1608; // @[Sbuffer.scala 134:17]
  wire  _GEN_3657 = line_mask_clean_valid_1 ? _GEN_2633 : _GEN_1609; // @[Sbuffer.scala 134:17]
  wire  _GEN_3658 = line_mask_clean_valid_1 ? _GEN_2634 : _GEN_1610; // @[Sbuffer.scala 134:17]
  wire  _GEN_3659 = line_mask_clean_valid_1 ? _GEN_2635 : _GEN_1611; // @[Sbuffer.scala 134:17]
  wire  _GEN_3660 = line_mask_clean_valid_1 ? _GEN_2636 : _GEN_1612; // @[Sbuffer.scala 134:17]
  wire  _GEN_3661 = line_mask_clean_valid_1 ? _GEN_2637 : _GEN_1613; // @[Sbuffer.scala 134:17]
  wire  _GEN_3662 = line_mask_clean_valid_1 ? _GEN_2638 : _GEN_1614; // @[Sbuffer.scala 134:17]
  wire  _GEN_3663 = line_mask_clean_valid_1 ? _GEN_2639 : _GEN_1615; // @[Sbuffer.scala 134:17]
  wire  _GEN_3664 = line_mask_clean_valid_1 ? _GEN_2640 : _GEN_1616; // @[Sbuffer.scala 134:17]
  wire  _GEN_3665 = line_mask_clean_valid_1 ? _GEN_2641 : _GEN_1617; // @[Sbuffer.scala 134:17]
  wire  _GEN_3666 = line_mask_clean_valid_1 ? _GEN_2642 : _GEN_1618; // @[Sbuffer.scala 134:17]
  wire  _GEN_3667 = line_mask_clean_valid_1 ? _GEN_2643 : _GEN_1619; // @[Sbuffer.scala 134:17]
  wire  _GEN_3668 = line_mask_clean_valid_1 ? _GEN_2644 : _GEN_1620; // @[Sbuffer.scala 134:17]
  wire  _GEN_3669 = line_mask_clean_valid_1 ? _GEN_2645 : _GEN_1621; // @[Sbuffer.scala 134:17]
  wire  _GEN_3670 = line_mask_clean_valid_1 ? _GEN_2646 : _GEN_1622; // @[Sbuffer.scala 134:17]
  wire  _GEN_3671 = line_mask_clean_valid_1 ? _GEN_2647 : _GEN_1623; // @[Sbuffer.scala 134:17]
  wire  _GEN_3672 = line_mask_clean_valid_1 ? _GEN_2648 : _GEN_1624; // @[Sbuffer.scala 134:17]
  wire  _GEN_3673 = line_mask_clean_valid_1 ? _GEN_2649 : _GEN_1625; // @[Sbuffer.scala 134:17]
  wire  _GEN_3674 = line_mask_clean_valid_1 ? _GEN_2650 : _GEN_1626; // @[Sbuffer.scala 134:17]
  wire  _GEN_3675 = line_mask_clean_valid_1 ? _GEN_2651 : _GEN_1627; // @[Sbuffer.scala 134:17]
  wire  _GEN_3676 = line_mask_clean_valid_1 ? _GEN_2652 : _GEN_1628; // @[Sbuffer.scala 134:17]
  wire  _GEN_3677 = line_mask_clean_valid_1 ? _GEN_2653 : _GEN_1629; // @[Sbuffer.scala 134:17]
  wire  _GEN_3678 = line_mask_clean_valid_1 ? _GEN_2654 : _GEN_1630; // @[Sbuffer.scala 134:17]
  wire  _GEN_3679 = line_mask_clean_valid_1 ? _GEN_2655 : _GEN_1631; // @[Sbuffer.scala 134:17]
  wire  _GEN_3680 = line_mask_clean_valid_1 ? _GEN_2656 : _GEN_1632; // @[Sbuffer.scala 134:17]
  wire  _GEN_3681 = line_mask_clean_valid_1 ? _GEN_2657 : _GEN_1633; // @[Sbuffer.scala 134:17]
  wire  _GEN_3682 = line_mask_clean_valid_1 ? _GEN_2658 : _GEN_1634; // @[Sbuffer.scala 134:17]
  wire  _GEN_3683 = line_mask_clean_valid_1 ? _GEN_2659 : _GEN_1635; // @[Sbuffer.scala 134:17]
  wire  _GEN_3684 = line_mask_clean_valid_1 ? _GEN_2660 : _GEN_1636; // @[Sbuffer.scala 134:17]
  wire  _GEN_3685 = line_mask_clean_valid_1 ? _GEN_2661 : _GEN_1637; // @[Sbuffer.scala 134:17]
  wire  _GEN_3686 = line_mask_clean_valid_1 ? _GEN_2662 : _GEN_1638; // @[Sbuffer.scala 134:17]
  wire  _GEN_3687 = line_mask_clean_valid_1 ? _GEN_2663 : _GEN_1639; // @[Sbuffer.scala 134:17]
  wire  _GEN_3688 = line_mask_clean_valid_1 ? _GEN_2664 : _GEN_1640; // @[Sbuffer.scala 134:17]
  wire  _GEN_3689 = line_mask_clean_valid_1 ? _GEN_2665 : _GEN_1641; // @[Sbuffer.scala 134:17]
  wire  _GEN_3690 = line_mask_clean_valid_1 ? _GEN_2666 : _GEN_1642; // @[Sbuffer.scala 134:17]
  wire  _GEN_3691 = line_mask_clean_valid_1 ? _GEN_2667 : _GEN_1643; // @[Sbuffer.scala 134:17]
  wire  _GEN_3692 = line_mask_clean_valid_1 ? _GEN_2668 : _GEN_1644; // @[Sbuffer.scala 134:17]
  wire  _GEN_3693 = line_mask_clean_valid_1 ? _GEN_2669 : _GEN_1645; // @[Sbuffer.scala 134:17]
  wire  _GEN_3694 = line_mask_clean_valid_1 ? _GEN_2670 : _GEN_1646; // @[Sbuffer.scala 134:17]
  wire  _GEN_3695 = line_mask_clean_valid_1 ? _GEN_2671 : _GEN_1647; // @[Sbuffer.scala 134:17]
  wire  _GEN_3696 = line_mask_clean_valid_1 ? _GEN_2672 : _GEN_1648; // @[Sbuffer.scala 134:17]
  wire  _GEN_3697 = line_mask_clean_valid_1 ? _GEN_2673 : _GEN_1649; // @[Sbuffer.scala 134:17]
  wire  _GEN_3698 = line_mask_clean_valid_1 ? _GEN_2674 : _GEN_1650; // @[Sbuffer.scala 134:17]
  wire  _GEN_3699 = line_mask_clean_valid_1 ? _GEN_2675 : _GEN_1651; // @[Sbuffer.scala 134:17]
  wire  _GEN_3700 = line_mask_clean_valid_1 ? _GEN_2676 : _GEN_1652; // @[Sbuffer.scala 134:17]
  wire  _GEN_3701 = line_mask_clean_valid_1 ? _GEN_2677 : _GEN_1653; // @[Sbuffer.scala 134:17]
  wire  _GEN_3702 = line_mask_clean_valid_1 ? _GEN_2678 : _GEN_1654; // @[Sbuffer.scala 134:17]
  wire  _GEN_3703 = line_mask_clean_valid_1 ? _GEN_2679 : _GEN_1655; // @[Sbuffer.scala 134:17]
  wire  _GEN_3704 = line_mask_clean_valid_1 ? _GEN_2680 : _GEN_1656; // @[Sbuffer.scala 134:17]
  wire  _GEN_3705 = line_mask_clean_valid_1 ? _GEN_2681 : _GEN_1657; // @[Sbuffer.scala 134:17]
  wire  _GEN_3706 = line_mask_clean_valid_1 ? _GEN_2682 : _GEN_1658; // @[Sbuffer.scala 134:17]
  wire  _GEN_3707 = line_mask_clean_valid_1 ? _GEN_2683 : _GEN_1659; // @[Sbuffer.scala 134:17]
  wire  _GEN_3708 = line_mask_clean_valid_1 ? _GEN_2684 : _GEN_1660; // @[Sbuffer.scala 134:17]
  wire  _GEN_3709 = line_mask_clean_valid_1 ? _GEN_2685 : _GEN_1661; // @[Sbuffer.scala 134:17]
  wire  _GEN_3710 = line_mask_clean_valid_1 ? _GEN_2686 : _GEN_1662; // @[Sbuffer.scala 134:17]
  wire  _GEN_3711 = line_mask_clean_valid_1 ? _GEN_2687 : _GEN_1663; // @[Sbuffer.scala 134:17]
  wire  _GEN_3712 = line_mask_clean_valid_1 ? _GEN_2688 : _GEN_1664; // @[Sbuffer.scala 134:17]
  wire  _GEN_3713 = line_mask_clean_valid_1 ? _GEN_2689 : _GEN_1665; // @[Sbuffer.scala 134:17]
  wire  _GEN_3714 = line_mask_clean_valid_1 ? _GEN_2690 : _GEN_1666; // @[Sbuffer.scala 134:17]
  wire  _GEN_3715 = line_mask_clean_valid_1 ? _GEN_2691 : _GEN_1667; // @[Sbuffer.scala 134:17]
  wire  _GEN_3716 = line_mask_clean_valid_1 ? _GEN_2692 : _GEN_1668; // @[Sbuffer.scala 134:17]
  wire  _GEN_3717 = line_mask_clean_valid_1 ? _GEN_2693 : _GEN_1669; // @[Sbuffer.scala 134:17]
  wire  _GEN_3718 = line_mask_clean_valid_1 ? _GEN_2694 : _GEN_1670; // @[Sbuffer.scala 134:17]
  wire  _GEN_3719 = line_mask_clean_valid_1 ? _GEN_2695 : _GEN_1671; // @[Sbuffer.scala 134:17]
  wire  _GEN_3720 = line_mask_clean_valid_1 ? _GEN_2696 : _GEN_1672; // @[Sbuffer.scala 134:17]
  wire  _GEN_3721 = line_mask_clean_valid_1 ? _GEN_2697 : _GEN_1673; // @[Sbuffer.scala 134:17]
  wire  _GEN_3722 = line_mask_clean_valid_1 ? _GEN_2698 : _GEN_1674; // @[Sbuffer.scala 134:17]
  wire  _GEN_3723 = line_mask_clean_valid_1 ? _GEN_2699 : _GEN_1675; // @[Sbuffer.scala 134:17]
  wire  _GEN_3724 = line_mask_clean_valid_1 ? _GEN_2700 : _GEN_1676; // @[Sbuffer.scala 134:17]
  wire  _GEN_3725 = line_mask_clean_valid_1 ? _GEN_2701 : _GEN_1677; // @[Sbuffer.scala 134:17]
  wire  _GEN_3726 = line_mask_clean_valid_1 ? _GEN_2702 : _GEN_1678; // @[Sbuffer.scala 134:17]
  wire  _GEN_3727 = line_mask_clean_valid_1 ? _GEN_2703 : _GEN_1679; // @[Sbuffer.scala 134:17]
  wire  _GEN_3728 = line_mask_clean_valid_1 ? _GEN_2704 : _GEN_1680; // @[Sbuffer.scala 134:17]
  wire  _GEN_3729 = line_mask_clean_valid_1 ? _GEN_2705 : _GEN_1681; // @[Sbuffer.scala 134:17]
  wire  _GEN_3730 = line_mask_clean_valid_1 ? _GEN_2706 : _GEN_1682; // @[Sbuffer.scala 134:17]
  wire  _GEN_3731 = line_mask_clean_valid_1 ? _GEN_2707 : _GEN_1683; // @[Sbuffer.scala 134:17]
  wire  _GEN_3732 = line_mask_clean_valid_1 ? _GEN_2708 : _GEN_1684; // @[Sbuffer.scala 134:17]
  wire  _GEN_3733 = line_mask_clean_valid_1 ? _GEN_2709 : _GEN_1685; // @[Sbuffer.scala 134:17]
  wire  _GEN_3734 = line_mask_clean_valid_1 ? _GEN_2710 : _GEN_1686; // @[Sbuffer.scala 134:17]
  wire  _GEN_3735 = line_mask_clean_valid_1 ? _GEN_2711 : _GEN_1687; // @[Sbuffer.scala 134:17]
  wire  _GEN_3736 = line_mask_clean_valid_1 ? _GEN_2712 : _GEN_1688; // @[Sbuffer.scala 134:17]
  wire  _GEN_3737 = line_mask_clean_valid_1 ? _GEN_2713 : _GEN_1689; // @[Sbuffer.scala 134:17]
  wire  _GEN_3738 = line_mask_clean_valid_1 ? _GEN_2714 : _GEN_1690; // @[Sbuffer.scala 134:17]
  wire  _GEN_3739 = line_mask_clean_valid_1 ? _GEN_2715 : _GEN_1691; // @[Sbuffer.scala 134:17]
  wire  _GEN_3740 = line_mask_clean_valid_1 ? _GEN_2716 : _GEN_1692; // @[Sbuffer.scala 134:17]
  wire  _GEN_3741 = line_mask_clean_valid_1 ? _GEN_2717 : _GEN_1693; // @[Sbuffer.scala 134:17]
  wire  _GEN_3742 = line_mask_clean_valid_1 ? _GEN_2718 : _GEN_1694; // @[Sbuffer.scala 134:17]
  wire  _GEN_3743 = line_mask_clean_valid_1 ? _GEN_2719 : _GEN_1695; // @[Sbuffer.scala 134:17]
  wire  _GEN_3744 = line_mask_clean_valid_1 ? _GEN_2720 : _GEN_1696; // @[Sbuffer.scala 134:17]
  wire  _GEN_3745 = line_mask_clean_valid_1 ? _GEN_2721 : _GEN_1697; // @[Sbuffer.scala 134:17]
  wire  _GEN_3746 = line_mask_clean_valid_1 ? _GEN_2722 : _GEN_1698; // @[Sbuffer.scala 134:17]
  wire  _GEN_3747 = line_mask_clean_valid_1 ? _GEN_2723 : _GEN_1699; // @[Sbuffer.scala 134:17]
  wire  _GEN_3748 = line_mask_clean_valid_1 ? _GEN_2724 : _GEN_1700; // @[Sbuffer.scala 134:17]
  wire  _GEN_3749 = line_mask_clean_valid_1 ? _GEN_2725 : _GEN_1701; // @[Sbuffer.scala 134:17]
  wire  _GEN_3750 = line_mask_clean_valid_1 ? _GEN_2726 : _GEN_1702; // @[Sbuffer.scala 134:17]
  wire  _GEN_3751 = line_mask_clean_valid_1 ? _GEN_2727 : _GEN_1703; // @[Sbuffer.scala 134:17]
  wire  _GEN_3752 = line_mask_clean_valid_1 ? _GEN_2728 : _GEN_1704; // @[Sbuffer.scala 134:17]
  wire  _GEN_3753 = line_mask_clean_valid_1 ? _GEN_2729 : _GEN_1705; // @[Sbuffer.scala 134:17]
  wire  _GEN_3754 = line_mask_clean_valid_1 ? _GEN_2730 : _GEN_1706; // @[Sbuffer.scala 134:17]
  wire  _GEN_3755 = line_mask_clean_valid_1 ? _GEN_2731 : _GEN_1707; // @[Sbuffer.scala 134:17]
  wire  _GEN_3756 = line_mask_clean_valid_1 ? _GEN_2732 : _GEN_1708; // @[Sbuffer.scala 134:17]
  wire  _GEN_3757 = line_mask_clean_valid_1 ? _GEN_2733 : _GEN_1709; // @[Sbuffer.scala 134:17]
  wire  _GEN_3758 = line_mask_clean_valid_1 ? _GEN_2734 : _GEN_1710; // @[Sbuffer.scala 134:17]
  wire  _GEN_3759 = line_mask_clean_valid_1 ? _GEN_2735 : _GEN_1711; // @[Sbuffer.scala 134:17]
  wire  _GEN_3760 = line_mask_clean_valid_1 ? _GEN_2736 : _GEN_1712; // @[Sbuffer.scala 134:17]
  wire  _GEN_3761 = line_mask_clean_valid_1 ? _GEN_2737 : _GEN_1713; // @[Sbuffer.scala 134:17]
  wire  _GEN_3762 = line_mask_clean_valid_1 ? _GEN_2738 : _GEN_1714; // @[Sbuffer.scala 134:17]
  wire  _GEN_3763 = line_mask_clean_valid_1 ? _GEN_2739 : _GEN_1715; // @[Sbuffer.scala 134:17]
  wire  _GEN_3764 = line_mask_clean_valid_1 ? _GEN_2740 : _GEN_1716; // @[Sbuffer.scala 134:17]
  wire  _GEN_3765 = line_mask_clean_valid_1 ? _GEN_2741 : _GEN_1717; // @[Sbuffer.scala 134:17]
  wire  _GEN_3766 = line_mask_clean_valid_1 ? _GEN_2742 : _GEN_1718; // @[Sbuffer.scala 134:17]
  wire  _GEN_3767 = line_mask_clean_valid_1 ? _GEN_2743 : _GEN_1719; // @[Sbuffer.scala 134:17]
  wire  _GEN_3768 = line_mask_clean_valid_1 ? _GEN_2744 : _GEN_1720; // @[Sbuffer.scala 134:17]
  wire  _GEN_3769 = line_mask_clean_valid_1 ? _GEN_2745 : _GEN_1721; // @[Sbuffer.scala 134:17]
  wire  _GEN_3770 = line_mask_clean_valid_1 ? _GEN_2746 : _GEN_1722; // @[Sbuffer.scala 134:17]
  wire  _GEN_3771 = line_mask_clean_valid_1 ? _GEN_2747 : _GEN_1723; // @[Sbuffer.scala 134:17]
  wire  _GEN_3772 = line_mask_clean_valid_1 ? _GEN_2748 : _GEN_1724; // @[Sbuffer.scala 134:17]
  wire  _GEN_3773 = line_mask_clean_valid_1 ? _GEN_2749 : _GEN_1725; // @[Sbuffer.scala 134:17]
  wire  _GEN_3774 = line_mask_clean_valid_1 ? _GEN_2750 : _GEN_1726; // @[Sbuffer.scala 134:17]
  wire  _GEN_3775 = line_mask_clean_valid_1 ? _GEN_2751 : _GEN_1727; // @[Sbuffer.scala 134:17]
  wire  _GEN_3776 = line_mask_clean_valid_1 ? _GEN_2752 : _GEN_1728; // @[Sbuffer.scala 134:17]
  wire  _GEN_3777 = line_mask_clean_valid_1 ? _GEN_2753 : _GEN_1729; // @[Sbuffer.scala 134:17]
  wire  _GEN_3778 = line_mask_clean_valid_1 ? _GEN_2754 : _GEN_1730; // @[Sbuffer.scala 134:17]
  wire  _GEN_3779 = line_mask_clean_valid_1 ? _GEN_2755 : _GEN_1731; // @[Sbuffer.scala 134:17]
  wire  _GEN_3780 = line_mask_clean_valid_1 ? _GEN_2756 : _GEN_1732; // @[Sbuffer.scala 134:17]
  wire  _GEN_3781 = line_mask_clean_valid_1 ? _GEN_2757 : _GEN_1733; // @[Sbuffer.scala 134:17]
  wire  _GEN_3782 = line_mask_clean_valid_1 ? _GEN_2758 : _GEN_1734; // @[Sbuffer.scala 134:17]
  wire  _GEN_3783 = line_mask_clean_valid_1 ? _GEN_2759 : _GEN_1735; // @[Sbuffer.scala 134:17]
  wire  _GEN_3784 = line_mask_clean_valid_1 ? _GEN_2760 : _GEN_1736; // @[Sbuffer.scala 134:17]
  wire  _GEN_3785 = line_mask_clean_valid_1 ? _GEN_2761 : _GEN_1737; // @[Sbuffer.scala 134:17]
  wire  _GEN_3786 = line_mask_clean_valid_1 ? _GEN_2762 : _GEN_1738; // @[Sbuffer.scala 134:17]
  wire  _GEN_3787 = line_mask_clean_valid_1 ? _GEN_2763 : _GEN_1739; // @[Sbuffer.scala 134:17]
  wire  _GEN_3788 = line_mask_clean_valid_1 ? _GEN_2764 : _GEN_1740; // @[Sbuffer.scala 134:17]
  wire  _GEN_3789 = line_mask_clean_valid_1 ? _GEN_2765 : _GEN_1741; // @[Sbuffer.scala 134:17]
  wire  _GEN_3790 = line_mask_clean_valid_1 ? _GEN_2766 : _GEN_1742; // @[Sbuffer.scala 134:17]
  wire  _GEN_3791 = line_mask_clean_valid_1 ? _GEN_2767 : _GEN_1743; // @[Sbuffer.scala 134:17]
  wire  _GEN_3792 = line_mask_clean_valid_1 ? _GEN_2768 : _GEN_1744; // @[Sbuffer.scala 134:17]
  wire  _GEN_3793 = line_mask_clean_valid_1 ? _GEN_2769 : _GEN_1745; // @[Sbuffer.scala 134:17]
  wire  _GEN_3794 = line_mask_clean_valid_1 ? _GEN_2770 : _GEN_1746; // @[Sbuffer.scala 134:17]
  wire  _GEN_3795 = line_mask_clean_valid_1 ? _GEN_2771 : _GEN_1747; // @[Sbuffer.scala 134:17]
  wire  _GEN_3796 = line_mask_clean_valid_1 ? _GEN_2772 : _GEN_1748; // @[Sbuffer.scala 134:17]
  wire  _GEN_3797 = line_mask_clean_valid_1 ? _GEN_2773 : _GEN_1749; // @[Sbuffer.scala 134:17]
  wire  _GEN_3798 = line_mask_clean_valid_1 ? _GEN_2774 : _GEN_1750; // @[Sbuffer.scala 134:17]
  wire  _GEN_3799 = line_mask_clean_valid_1 ? _GEN_2775 : _GEN_1751; // @[Sbuffer.scala 134:17]
  wire  _GEN_3800 = line_mask_clean_valid_1 ? _GEN_2776 : _GEN_1752; // @[Sbuffer.scala 134:17]
  wire  _GEN_3801 = line_mask_clean_valid_1 ? _GEN_2777 : _GEN_1753; // @[Sbuffer.scala 134:17]
  wire  _GEN_3802 = line_mask_clean_valid_1 ? _GEN_2778 : _GEN_1754; // @[Sbuffer.scala 134:17]
  wire  _GEN_3803 = line_mask_clean_valid_1 ? _GEN_2779 : _GEN_1755; // @[Sbuffer.scala 134:17]
  wire  _GEN_3804 = line_mask_clean_valid_1 ? _GEN_2780 : _GEN_1756; // @[Sbuffer.scala 134:17]
  wire  _GEN_3805 = line_mask_clean_valid_1 ? _GEN_2781 : _GEN_1757; // @[Sbuffer.scala 134:17]
  wire  _GEN_3806 = line_mask_clean_valid_1 ? _GEN_2782 : _GEN_1758; // @[Sbuffer.scala 134:17]
  wire  _GEN_3807 = line_mask_clean_valid_1 ? _GEN_2783 : _GEN_1759; // @[Sbuffer.scala 134:17]
  wire  _GEN_3808 = line_mask_clean_valid_1 ? _GEN_2784 : _GEN_1760; // @[Sbuffer.scala 134:17]
  wire  _GEN_3809 = line_mask_clean_valid_1 ? _GEN_2785 : _GEN_1761; // @[Sbuffer.scala 134:17]
  wire  _GEN_3810 = line_mask_clean_valid_1 ? _GEN_2786 : _GEN_1762; // @[Sbuffer.scala 134:17]
  wire  _GEN_3811 = line_mask_clean_valid_1 ? _GEN_2787 : _GEN_1763; // @[Sbuffer.scala 134:17]
  wire  _GEN_3812 = line_mask_clean_valid_1 ? _GEN_2788 : _GEN_1764; // @[Sbuffer.scala 134:17]
  wire  _GEN_3813 = line_mask_clean_valid_1 ? _GEN_2789 : _GEN_1765; // @[Sbuffer.scala 134:17]
  wire  _GEN_3814 = line_mask_clean_valid_1 ? _GEN_2790 : _GEN_1766; // @[Sbuffer.scala 134:17]
  wire  _GEN_3815 = line_mask_clean_valid_1 ? _GEN_2791 : _GEN_1767; // @[Sbuffer.scala 134:17]
  wire  _GEN_3816 = line_mask_clean_valid_1 ? _GEN_2792 : _GEN_1768; // @[Sbuffer.scala 134:17]
  wire  _GEN_3817 = line_mask_clean_valid_1 ? _GEN_2793 : _GEN_1769; // @[Sbuffer.scala 134:17]
  wire  _GEN_3818 = line_mask_clean_valid_1 ? _GEN_2794 : _GEN_1770; // @[Sbuffer.scala 134:17]
  wire  _GEN_3819 = line_mask_clean_valid_1 ? _GEN_2795 : _GEN_1771; // @[Sbuffer.scala 134:17]
  wire  _GEN_3820 = line_mask_clean_valid_1 ? _GEN_2796 : _GEN_1772; // @[Sbuffer.scala 134:17]
  wire  _GEN_3821 = line_mask_clean_valid_1 ? _GEN_2797 : _GEN_1773; // @[Sbuffer.scala 134:17]
  wire  _GEN_3822 = line_mask_clean_valid_1 ? _GEN_2798 : _GEN_1774; // @[Sbuffer.scala 134:17]
  wire  _GEN_3823 = line_mask_clean_valid_1 ? _GEN_2799 : _GEN_1775; // @[Sbuffer.scala 134:17]
  wire  _GEN_3824 = line_mask_clean_valid_1 ? _GEN_2800 : _GEN_1776; // @[Sbuffer.scala 134:17]
  wire  _GEN_3825 = line_mask_clean_valid_1 ? _GEN_2801 : _GEN_1777; // @[Sbuffer.scala 134:17]
  wire  _GEN_3826 = line_mask_clean_valid_1 ? _GEN_2802 : _GEN_1778; // @[Sbuffer.scala 134:17]
  wire  _GEN_3827 = line_mask_clean_valid_1 ? _GEN_2803 : _GEN_1779; // @[Sbuffer.scala 134:17]
  wire  _GEN_3828 = line_mask_clean_valid_1 ? _GEN_2804 : _GEN_1780; // @[Sbuffer.scala 134:17]
  wire  _GEN_3829 = line_mask_clean_valid_1 ? _GEN_2805 : _GEN_1781; // @[Sbuffer.scala 134:17]
  wire  _GEN_3830 = line_mask_clean_valid_1 ? _GEN_2806 : _GEN_1782; // @[Sbuffer.scala 134:17]
  wire  _GEN_3831 = line_mask_clean_valid_1 ? _GEN_2807 : _GEN_1783; // @[Sbuffer.scala 134:17]
  wire  _GEN_3832 = line_mask_clean_valid_1 ? _GEN_2808 : _GEN_1784; // @[Sbuffer.scala 134:17]
  wire  _GEN_3833 = line_mask_clean_valid_1 ? _GEN_2809 : _GEN_1785; // @[Sbuffer.scala 134:17]
  wire  _GEN_3834 = line_mask_clean_valid_1 ? _GEN_2810 : _GEN_1786; // @[Sbuffer.scala 134:17]
  wire  _GEN_3835 = line_mask_clean_valid_1 ? _GEN_2811 : _GEN_1787; // @[Sbuffer.scala 134:17]
  wire  _GEN_3836 = line_mask_clean_valid_1 ? _GEN_2812 : _GEN_1788; // @[Sbuffer.scala 134:17]
  wire  _GEN_3837 = line_mask_clean_valid_1 ? _GEN_2813 : _GEN_1789; // @[Sbuffer.scala 134:17]
  wire  _GEN_3838 = line_mask_clean_valid_1 ? _GEN_2814 : _GEN_1790; // @[Sbuffer.scala 134:17]
  wire  _GEN_3839 = line_mask_clean_valid_1 ? _GEN_2815 : _GEN_1791; // @[Sbuffer.scala 134:17]
  wire  _GEN_3840 = line_mask_clean_valid_1 ? _GEN_2816 : _GEN_1792; // @[Sbuffer.scala 134:17]
  wire  _GEN_3841 = line_mask_clean_valid_1 ? _GEN_2817 : _GEN_1793; // @[Sbuffer.scala 134:17]
  wire  _GEN_3842 = line_mask_clean_valid_1 ? _GEN_2818 : _GEN_1794; // @[Sbuffer.scala 134:17]
  wire  _GEN_3843 = line_mask_clean_valid_1 ? _GEN_2819 : _GEN_1795; // @[Sbuffer.scala 134:17]
  wire  _GEN_3844 = line_mask_clean_valid_1 ? _GEN_2820 : _GEN_1796; // @[Sbuffer.scala 134:17]
  wire  _GEN_3845 = line_mask_clean_valid_1 ? _GEN_2821 : _GEN_1797; // @[Sbuffer.scala 134:17]
  wire  _GEN_3846 = line_mask_clean_valid_1 ? _GEN_2822 : _GEN_1798; // @[Sbuffer.scala 134:17]
  wire  _GEN_3847 = line_mask_clean_valid_1 ? _GEN_2823 : _GEN_1799; // @[Sbuffer.scala 134:17]
  wire  _GEN_3848 = line_mask_clean_valid_1 ? _GEN_2824 : _GEN_1800; // @[Sbuffer.scala 134:17]
  wire  _GEN_3849 = line_mask_clean_valid_1 ? _GEN_2825 : _GEN_1801; // @[Sbuffer.scala 134:17]
  wire  _GEN_3850 = line_mask_clean_valid_1 ? _GEN_2826 : _GEN_1802; // @[Sbuffer.scala 134:17]
  wire  _GEN_3851 = line_mask_clean_valid_1 ? _GEN_2827 : _GEN_1803; // @[Sbuffer.scala 134:17]
  wire  _GEN_3852 = line_mask_clean_valid_1 ? _GEN_2828 : _GEN_1804; // @[Sbuffer.scala 134:17]
  wire  _GEN_3853 = line_mask_clean_valid_1 ? _GEN_2829 : _GEN_1805; // @[Sbuffer.scala 134:17]
  wire  _GEN_3854 = line_mask_clean_valid_1 ? _GEN_2830 : _GEN_1806; // @[Sbuffer.scala 134:17]
  wire  _GEN_3855 = line_mask_clean_valid_1 ? _GEN_2831 : _GEN_1807; // @[Sbuffer.scala 134:17]
  wire  _GEN_3856 = line_mask_clean_valid_1 ? _GEN_2832 : _GEN_1808; // @[Sbuffer.scala 134:17]
  wire  _GEN_3857 = line_mask_clean_valid_1 ? _GEN_2833 : _GEN_1809; // @[Sbuffer.scala 134:17]
  wire  _GEN_3858 = line_mask_clean_valid_1 ? _GEN_2834 : _GEN_1810; // @[Sbuffer.scala 134:17]
  wire  _GEN_3859 = line_mask_clean_valid_1 ? _GEN_2835 : _GEN_1811; // @[Sbuffer.scala 134:17]
  wire  _GEN_3860 = line_mask_clean_valid_1 ? _GEN_2836 : _GEN_1812; // @[Sbuffer.scala 134:17]
  wire  _GEN_3861 = line_mask_clean_valid_1 ? _GEN_2837 : _GEN_1813; // @[Sbuffer.scala 134:17]
  wire  _GEN_3862 = line_mask_clean_valid_1 ? _GEN_2838 : _GEN_1814; // @[Sbuffer.scala 134:17]
  wire  _GEN_3863 = line_mask_clean_valid_1 ? _GEN_2839 : _GEN_1815; // @[Sbuffer.scala 134:17]
  wire  _GEN_3864 = line_mask_clean_valid_1 ? _GEN_2840 : _GEN_1816; // @[Sbuffer.scala 134:17]
  wire  _GEN_3865 = line_mask_clean_valid_1 ? _GEN_2841 : _GEN_1817; // @[Sbuffer.scala 134:17]
  wire  _GEN_3866 = line_mask_clean_valid_1 ? _GEN_2842 : _GEN_1818; // @[Sbuffer.scala 134:17]
  wire  _GEN_3867 = line_mask_clean_valid_1 ? _GEN_2843 : _GEN_1819; // @[Sbuffer.scala 134:17]
  wire  _GEN_3868 = line_mask_clean_valid_1 ? _GEN_2844 : _GEN_1820; // @[Sbuffer.scala 134:17]
  wire  _GEN_3869 = line_mask_clean_valid_1 ? _GEN_2845 : _GEN_1821; // @[Sbuffer.scala 134:17]
  wire  _GEN_3870 = line_mask_clean_valid_1 ? _GEN_2846 : _GEN_1822; // @[Sbuffer.scala 134:17]
  wire  _GEN_3871 = line_mask_clean_valid_1 ? _GEN_2847 : _GEN_1823; // @[Sbuffer.scala 134:17]
  wire  _GEN_3872 = line_mask_clean_valid_1 ? _GEN_2848 : _GEN_1824; // @[Sbuffer.scala 134:17]
  wire  _GEN_3873 = line_mask_clean_valid_1 ? _GEN_2849 : _GEN_1825; // @[Sbuffer.scala 134:17]
  wire  _GEN_3874 = line_mask_clean_valid_1 ? _GEN_2850 : _GEN_1826; // @[Sbuffer.scala 134:17]
  wire  _GEN_3875 = line_mask_clean_valid_1 ? _GEN_2851 : _GEN_1827; // @[Sbuffer.scala 134:17]
  wire  _GEN_3876 = line_mask_clean_valid_1 ? _GEN_2852 : _GEN_1828; // @[Sbuffer.scala 134:17]
  wire  _GEN_3877 = line_mask_clean_valid_1 ? _GEN_2853 : _GEN_1829; // @[Sbuffer.scala 134:17]
  wire  _GEN_3878 = line_mask_clean_valid_1 ? _GEN_2854 : _GEN_1830; // @[Sbuffer.scala 134:17]
  wire  _GEN_3879 = line_mask_clean_valid_1 ? _GEN_2855 : _GEN_1831; // @[Sbuffer.scala 134:17]
  wire  _GEN_3880 = line_mask_clean_valid_1 ? _GEN_2856 : _GEN_1832; // @[Sbuffer.scala 134:17]
  wire  _GEN_3881 = line_mask_clean_valid_1 ? _GEN_2857 : _GEN_1833; // @[Sbuffer.scala 134:17]
  wire  _GEN_3882 = line_mask_clean_valid_1 ? _GEN_2858 : _GEN_1834; // @[Sbuffer.scala 134:17]
  wire  _GEN_3883 = line_mask_clean_valid_1 ? _GEN_2859 : _GEN_1835; // @[Sbuffer.scala 134:17]
  wire  _GEN_3884 = line_mask_clean_valid_1 ? _GEN_2860 : _GEN_1836; // @[Sbuffer.scala 134:17]
  wire  _GEN_3885 = line_mask_clean_valid_1 ? _GEN_2861 : _GEN_1837; // @[Sbuffer.scala 134:17]
  wire  _GEN_3886 = line_mask_clean_valid_1 ? _GEN_2862 : _GEN_1838; // @[Sbuffer.scala 134:17]
  wire  _GEN_3887 = line_mask_clean_valid_1 ? _GEN_2863 : _GEN_1839; // @[Sbuffer.scala 134:17]
  wire  _GEN_3888 = line_mask_clean_valid_1 ? _GEN_2864 : _GEN_1840; // @[Sbuffer.scala 134:17]
  wire  _GEN_3889 = line_mask_clean_valid_1 ? _GEN_2865 : _GEN_1841; // @[Sbuffer.scala 134:17]
  wire  _GEN_3890 = line_mask_clean_valid_1 ? _GEN_2866 : _GEN_1842; // @[Sbuffer.scala 134:17]
  wire  _GEN_3891 = line_mask_clean_valid_1 ? _GEN_2867 : _GEN_1843; // @[Sbuffer.scala 134:17]
  wire  _GEN_3892 = line_mask_clean_valid_1 ? _GEN_2868 : _GEN_1844; // @[Sbuffer.scala 134:17]
  wire  _GEN_3893 = line_mask_clean_valid_1 ? _GEN_2869 : _GEN_1845; // @[Sbuffer.scala 134:17]
  wire  _GEN_3894 = line_mask_clean_valid_1 ? _GEN_2870 : _GEN_1846; // @[Sbuffer.scala 134:17]
  wire  _GEN_3895 = line_mask_clean_valid_1 ? _GEN_2871 : _GEN_1847; // @[Sbuffer.scala 134:17]
  wire  _GEN_3896 = line_mask_clean_valid_1 ? _GEN_2872 : _GEN_1848; // @[Sbuffer.scala 134:17]
  wire  _GEN_3897 = line_mask_clean_valid_1 ? _GEN_2873 : _GEN_1849; // @[Sbuffer.scala 134:17]
  wire  _GEN_3898 = line_mask_clean_valid_1 ? _GEN_2874 : _GEN_1850; // @[Sbuffer.scala 134:17]
  wire  _GEN_3899 = line_mask_clean_valid_1 ? _GEN_2875 : _GEN_1851; // @[Sbuffer.scala 134:17]
  wire  _GEN_3900 = line_mask_clean_valid_1 ? _GEN_2876 : _GEN_1852; // @[Sbuffer.scala 134:17]
  wire  _GEN_3901 = line_mask_clean_valid_1 ? _GEN_2877 : _GEN_1853; // @[Sbuffer.scala 134:17]
  wire  _GEN_3902 = line_mask_clean_valid_1 ? _GEN_2878 : _GEN_1854; // @[Sbuffer.scala 134:17]
  wire  _GEN_3903 = line_mask_clean_valid_1 ? _GEN_2879 : _GEN_1855; // @[Sbuffer.scala 134:17]
  wire  _GEN_3904 = line_mask_clean_valid_1 ? _GEN_2880 : _GEN_1856; // @[Sbuffer.scala 134:17]
  wire  _GEN_3905 = line_mask_clean_valid_1 ? _GEN_2881 : _GEN_1857; // @[Sbuffer.scala 134:17]
  wire  _GEN_3906 = line_mask_clean_valid_1 ? _GEN_2882 : _GEN_1858; // @[Sbuffer.scala 134:17]
  wire  _GEN_3907 = line_mask_clean_valid_1 ? _GEN_2883 : _GEN_1859; // @[Sbuffer.scala 134:17]
  wire  _GEN_3908 = line_mask_clean_valid_1 ? _GEN_2884 : _GEN_1860; // @[Sbuffer.scala 134:17]
  wire  _GEN_3909 = line_mask_clean_valid_1 ? _GEN_2885 : _GEN_1861; // @[Sbuffer.scala 134:17]
  wire  _GEN_3910 = line_mask_clean_valid_1 ? _GEN_2886 : _GEN_1862; // @[Sbuffer.scala 134:17]
  wire  _GEN_3911 = line_mask_clean_valid_1 ? _GEN_2887 : _GEN_1863; // @[Sbuffer.scala 134:17]
  wire  _GEN_3912 = line_mask_clean_valid_1 ? _GEN_2888 : _GEN_1864; // @[Sbuffer.scala 134:17]
  wire  _GEN_3913 = line_mask_clean_valid_1 ? _GEN_2889 : _GEN_1865; // @[Sbuffer.scala 134:17]
  wire  _GEN_3914 = line_mask_clean_valid_1 ? _GEN_2890 : _GEN_1866; // @[Sbuffer.scala 134:17]
  wire  _GEN_3915 = line_mask_clean_valid_1 ? _GEN_2891 : _GEN_1867; // @[Sbuffer.scala 134:17]
  wire  _GEN_3916 = line_mask_clean_valid_1 ? _GEN_2892 : _GEN_1868; // @[Sbuffer.scala 134:17]
  wire  _GEN_3917 = line_mask_clean_valid_1 ? _GEN_2893 : _GEN_1869; // @[Sbuffer.scala 134:17]
  wire  _GEN_3918 = line_mask_clean_valid_1 ? _GEN_2894 : _GEN_1870; // @[Sbuffer.scala 134:17]
  wire  _GEN_3919 = line_mask_clean_valid_1 ? _GEN_2895 : _GEN_1871; // @[Sbuffer.scala 134:17]
  wire  _GEN_3920 = line_mask_clean_valid_1 ? _GEN_2896 : _GEN_1872; // @[Sbuffer.scala 134:17]
  wire  _GEN_3921 = line_mask_clean_valid_1 ? _GEN_2897 : _GEN_1873; // @[Sbuffer.scala 134:17]
  wire  _GEN_3922 = line_mask_clean_valid_1 ? _GEN_2898 : _GEN_1874; // @[Sbuffer.scala 134:17]
  wire  _GEN_3923 = line_mask_clean_valid_1 ? _GEN_2899 : _GEN_1875; // @[Sbuffer.scala 134:17]
  wire  _GEN_3924 = line_mask_clean_valid_1 ? _GEN_2900 : _GEN_1876; // @[Sbuffer.scala 134:17]
  wire  _GEN_3925 = line_mask_clean_valid_1 ? _GEN_2901 : _GEN_1877; // @[Sbuffer.scala 134:17]
  wire  _GEN_3926 = line_mask_clean_valid_1 ? _GEN_2902 : _GEN_1878; // @[Sbuffer.scala 134:17]
  wire  _GEN_3927 = line_mask_clean_valid_1 ? _GEN_2903 : _GEN_1879; // @[Sbuffer.scala 134:17]
  wire  _GEN_3928 = line_mask_clean_valid_1 ? _GEN_2904 : _GEN_1880; // @[Sbuffer.scala 134:17]
  wire  _GEN_3929 = line_mask_clean_valid_1 ? _GEN_2905 : _GEN_1881; // @[Sbuffer.scala 134:17]
  wire  _GEN_3930 = line_mask_clean_valid_1 ? _GEN_2906 : _GEN_1882; // @[Sbuffer.scala 134:17]
  wire  _GEN_3931 = line_mask_clean_valid_1 ? _GEN_2907 : _GEN_1883; // @[Sbuffer.scala 134:17]
  wire  _GEN_3932 = line_mask_clean_valid_1 ? _GEN_2908 : _GEN_1884; // @[Sbuffer.scala 134:17]
  wire  _GEN_3933 = line_mask_clean_valid_1 ? _GEN_2909 : _GEN_1885; // @[Sbuffer.scala 134:17]
  wire  _GEN_3934 = line_mask_clean_valid_1 ? _GEN_2910 : _GEN_1886; // @[Sbuffer.scala 134:17]
  wire  _GEN_3935 = line_mask_clean_valid_1 ? _GEN_2911 : _GEN_1887; // @[Sbuffer.scala 134:17]
  wire  _GEN_3936 = line_mask_clean_valid_1 ? _GEN_2912 : _GEN_1888; // @[Sbuffer.scala 134:17]
  wire  _GEN_3937 = line_mask_clean_valid_1 ? _GEN_2913 : _GEN_1889; // @[Sbuffer.scala 134:17]
  wire  _GEN_3938 = line_mask_clean_valid_1 ? _GEN_2914 : _GEN_1890; // @[Sbuffer.scala 134:17]
  wire  _GEN_3939 = line_mask_clean_valid_1 ? _GEN_2915 : _GEN_1891; // @[Sbuffer.scala 134:17]
  wire  _GEN_3940 = line_mask_clean_valid_1 ? _GEN_2916 : _GEN_1892; // @[Sbuffer.scala 134:17]
  wire  _GEN_3941 = line_mask_clean_valid_1 ? _GEN_2917 : _GEN_1893; // @[Sbuffer.scala 134:17]
  wire  _GEN_3942 = line_mask_clean_valid_1 ? _GEN_2918 : _GEN_1894; // @[Sbuffer.scala 134:17]
  wire  _GEN_3943 = line_mask_clean_valid_1 ? _GEN_2919 : _GEN_1895; // @[Sbuffer.scala 134:17]
  wire  _GEN_3944 = line_mask_clean_valid_1 ? _GEN_2920 : _GEN_1896; // @[Sbuffer.scala 134:17]
  wire  _GEN_3945 = line_mask_clean_valid_1 ? _GEN_2921 : _GEN_1897; // @[Sbuffer.scala 134:17]
  wire  _GEN_3946 = line_mask_clean_valid_1 ? _GEN_2922 : _GEN_1898; // @[Sbuffer.scala 134:17]
  wire  _GEN_3947 = line_mask_clean_valid_1 ? _GEN_2923 : _GEN_1899; // @[Sbuffer.scala 134:17]
  wire  _GEN_3948 = line_mask_clean_valid_1 ? _GEN_2924 : _GEN_1900; // @[Sbuffer.scala 134:17]
  wire  _GEN_3949 = line_mask_clean_valid_1 ? _GEN_2925 : _GEN_1901; // @[Sbuffer.scala 134:17]
  wire  _GEN_3950 = line_mask_clean_valid_1 ? _GEN_2926 : _GEN_1902; // @[Sbuffer.scala 134:17]
  wire  _GEN_3951 = line_mask_clean_valid_1 ? _GEN_2927 : _GEN_1903; // @[Sbuffer.scala 134:17]
  wire  _GEN_3952 = line_mask_clean_valid_1 ? _GEN_2928 : _GEN_1904; // @[Sbuffer.scala 134:17]
  wire  _GEN_3953 = line_mask_clean_valid_1 ? _GEN_2929 : _GEN_1905; // @[Sbuffer.scala 134:17]
  wire  _GEN_3954 = line_mask_clean_valid_1 ? _GEN_2930 : _GEN_1906; // @[Sbuffer.scala 134:17]
  wire  _GEN_3955 = line_mask_clean_valid_1 ? _GEN_2931 : _GEN_1907; // @[Sbuffer.scala 134:17]
  wire  _GEN_3956 = line_mask_clean_valid_1 ? _GEN_2932 : _GEN_1908; // @[Sbuffer.scala 134:17]
  wire  _GEN_3957 = line_mask_clean_valid_1 ? _GEN_2933 : _GEN_1909; // @[Sbuffer.scala 134:17]
  wire  _GEN_3958 = line_mask_clean_valid_1 ? _GEN_2934 : _GEN_1910; // @[Sbuffer.scala 134:17]
  wire  _GEN_3959 = line_mask_clean_valid_1 ? _GEN_2935 : _GEN_1911; // @[Sbuffer.scala 134:17]
  wire  _GEN_3960 = line_mask_clean_valid_1 ? _GEN_2936 : _GEN_1912; // @[Sbuffer.scala 134:17]
  wire  _GEN_3961 = line_mask_clean_valid_1 ? _GEN_2937 : _GEN_1913; // @[Sbuffer.scala 134:17]
  wire  _GEN_3962 = line_mask_clean_valid_1 ? _GEN_2938 : _GEN_1914; // @[Sbuffer.scala 134:17]
  wire  _GEN_3963 = line_mask_clean_valid_1 ? _GEN_2939 : _GEN_1915; // @[Sbuffer.scala 134:17]
  wire  _GEN_3964 = line_mask_clean_valid_1 ? _GEN_2940 : _GEN_1916; // @[Sbuffer.scala 134:17]
  wire  _GEN_3965 = line_mask_clean_valid_1 ? _GEN_2941 : _GEN_1917; // @[Sbuffer.scala 134:17]
  wire  _GEN_3966 = line_mask_clean_valid_1 ? _GEN_2942 : _GEN_1918; // @[Sbuffer.scala 134:17]
  wire  _GEN_3967 = line_mask_clean_valid_1 ? _GEN_2943 : _GEN_1919; // @[Sbuffer.scala 134:17]
  wire  _GEN_3968 = line_mask_clean_valid_1 ? _GEN_2944 : _GEN_1920; // @[Sbuffer.scala 134:17]
  wire  _GEN_3969 = line_mask_clean_valid_1 ? _GEN_2945 : _GEN_1921; // @[Sbuffer.scala 134:17]
  wire  _GEN_3970 = line_mask_clean_valid_1 ? _GEN_2946 : _GEN_1922; // @[Sbuffer.scala 134:17]
  wire  _GEN_3971 = line_mask_clean_valid_1 ? _GEN_2947 : _GEN_1923; // @[Sbuffer.scala 134:17]
  wire  _GEN_3972 = line_mask_clean_valid_1 ? _GEN_2948 : _GEN_1924; // @[Sbuffer.scala 134:17]
  wire  _GEN_3973 = line_mask_clean_valid_1 ? _GEN_2949 : _GEN_1925; // @[Sbuffer.scala 134:17]
  wire  _GEN_3974 = line_mask_clean_valid_1 ? _GEN_2950 : _GEN_1926; // @[Sbuffer.scala 134:17]
  wire  _GEN_3975 = line_mask_clean_valid_1 ? _GEN_2951 : _GEN_1927; // @[Sbuffer.scala 134:17]
  wire  _GEN_3976 = line_mask_clean_valid_1 ? _GEN_2952 : _GEN_1928; // @[Sbuffer.scala 134:17]
  wire  _GEN_3977 = line_mask_clean_valid_1 ? _GEN_2953 : _GEN_1929; // @[Sbuffer.scala 134:17]
  wire  _GEN_3978 = line_mask_clean_valid_1 ? _GEN_2954 : _GEN_1930; // @[Sbuffer.scala 134:17]
  wire  _GEN_3979 = line_mask_clean_valid_1 ? _GEN_2955 : _GEN_1931; // @[Sbuffer.scala 134:17]
  wire  _GEN_3980 = line_mask_clean_valid_1 ? _GEN_2956 : _GEN_1932; // @[Sbuffer.scala 134:17]
  wire  _GEN_3981 = line_mask_clean_valid_1 ? _GEN_2957 : _GEN_1933; // @[Sbuffer.scala 134:17]
  wire  _GEN_3982 = line_mask_clean_valid_1 ? _GEN_2958 : _GEN_1934; // @[Sbuffer.scala 134:17]
  wire  _GEN_3983 = line_mask_clean_valid_1 ? _GEN_2959 : _GEN_1935; // @[Sbuffer.scala 134:17]
  wire  _GEN_3984 = line_mask_clean_valid_1 ? _GEN_2960 : _GEN_1936; // @[Sbuffer.scala 134:17]
  wire  _GEN_3985 = line_mask_clean_valid_1 ? _GEN_2961 : _GEN_1937; // @[Sbuffer.scala 134:17]
  wire  _GEN_3986 = line_mask_clean_valid_1 ? _GEN_2962 : _GEN_1938; // @[Sbuffer.scala 134:17]
  wire  _GEN_3987 = line_mask_clean_valid_1 ? _GEN_2963 : _GEN_1939; // @[Sbuffer.scala 134:17]
  wire  _GEN_3988 = line_mask_clean_valid_1 ? _GEN_2964 : _GEN_1940; // @[Sbuffer.scala 134:17]
  wire  _GEN_3989 = line_mask_clean_valid_1 ? _GEN_2965 : _GEN_1941; // @[Sbuffer.scala 134:17]
  wire  _GEN_3990 = line_mask_clean_valid_1 ? _GEN_2966 : _GEN_1942; // @[Sbuffer.scala 134:17]
  wire  _GEN_3991 = line_mask_clean_valid_1 ? _GEN_2967 : _GEN_1943; // @[Sbuffer.scala 134:17]
  wire  _GEN_3992 = line_mask_clean_valid_1 ? _GEN_2968 : _GEN_1944; // @[Sbuffer.scala 134:17]
  wire  _GEN_3993 = line_mask_clean_valid_1 ? _GEN_2969 : _GEN_1945; // @[Sbuffer.scala 134:17]
  wire  _GEN_3994 = line_mask_clean_valid_1 ? _GEN_2970 : _GEN_1946; // @[Sbuffer.scala 134:17]
  wire  _GEN_3995 = line_mask_clean_valid_1 ? _GEN_2971 : _GEN_1947; // @[Sbuffer.scala 134:17]
  wire  _GEN_3996 = line_mask_clean_valid_1 ? _GEN_2972 : _GEN_1948; // @[Sbuffer.scala 134:17]
  wire  _GEN_3997 = line_mask_clean_valid_1 ? _GEN_2973 : _GEN_1949; // @[Sbuffer.scala 134:17]
  wire  _GEN_3998 = line_mask_clean_valid_1 ? _GEN_2974 : _GEN_1950; // @[Sbuffer.scala 134:17]
  wire  _GEN_3999 = line_mask_clean_valid_1 ? _GEN_2975 : _GEN_1951; // @[Sbuffer.scala 134:17]
  wire  _GEN_4000 = line_mask_clean_valid_1 ? _GEN_2976 : _GEN_1952; // @[Sbuffer.scala 134:17]
  wire  _GEN_4001 = line_mask_clean_valid_1 ? _GEN_2977 : _GEN_1953; // @[Sbuffer.scala 134:17]
  wire  _GEN_4002 = line_mask_clean_valid_1 ? _GEN_2978 : _GEN_1954; // @[Sbuffer.scala 134:17]
  wire  _GEN_4003 = line_mask_clean_valid_1 ? _GEN_2979 : _GEN_1955; // @[Sbuffer.scala 134:17]
  wire  _GEN_4004 = line_mask_clean_valid_1 ? _GEN_2980 : _GEN_1956; // @[Sbuffer.scala 134:17]
  wire  _GEN_4005 = line_mask_clean_valid_1 ? _GEN_2981 : _GEN_1957; // @[Sbuffer.scala 134:17]
  wire  _GEN_4006 = line_mask_clean_valid_1 ? _GEN_2982 : _GEN_1958; // @[Sbuffer.scala 134:17]
  wire  _GEN_4007 = line_mask_clean_valid_1 ? _GEN_2983 : _GEN_1959; // @[Sbuffer.scala 134:17]
  wire  _GEN_4008 = line_mask_clean_valid_1 ? _GEN_2984 : _GEN_1960; // @[Sbuffer.scala 134:17]
  wire  _GEN_4009 = line_mask_clean_valid_1 ? _GEN_2985 : _GEN_1961; // @[Sbuffer.scala 134:17]
  wire  _GEN_4010 = line_mask_clean_valid_1 ? _GEN_2986 : _GEN_1962; // @[Sbuffer.scala 134:17]
  wire  _GEN_4011 = line_mask_clean_valid_1 ? _GEN_2987 : _GEN_1963; // @[Sbuffer.scala 134:17]
  wire  _GEN_4012 = line_mask_clean_valid_1 ? _GEN_2988 : _GEN_1964; // @[Sbuffer.scala 134:17]
  wire  _GEN_4013 = line_mask_clean_valid_1 ? _GEN_2989 : _GEN_1965; // @[Sbuffer.scala 134:17]
  wire  _GEN_4014 = line_mask_clean_valid_1 ? _GEN_2990 : _GEN_1966; // @[Sbuffer.scala 134:17]
  wire  _GEN_4015 = line_mask_clean_valid_1 ? _GEN_2991 : _GEN_1967; // @[Sbuffer.scala 134:17]
  wire  _GEN_4016 = line_mask_clean_valid_1 ? _GEN_2992 : _GEN_1968; // @[Sbuffer.scala 134:17]
  wire  _GEN_4017 = line_mask_clean_valid_1 ? _GEN_2993 : _GEN_1969; // @[Sbuffer.scala 134:17]
  wire  _GEN_4018 = line_mask_clean_valid_1 ? _GEN_2994 : _GEN_1970; // @[Sbuffer.scala 134:17]
  wire  _GEN_4019 = line_mask_clean_valid_1 ? _GEN_2995 : _GEN_1971; // @[Sbuffer.scala 134:17]
  wire  _GEN_4020 = line_mask_clean_valid_1 ? _GEN_2996 : _GEN_1972; // @[Sbuffer.scala 134:17]
  wire  _GEN_4021 = line_mask_clean_valid_1 ? _GEN_2997 : _GEN_1973; // @[Sbuffer.scala 134:17]
  wire  _GEN_4022 = line_mask_clean_valid_1 ? _GEN_2998 : _GEN_1974; // @[Sbuffer.scala 134:17]
  wire  _GEN_4023 = line_mask_clean_valid_1 ? _GEN_2999 : _GEN_1975; // @[Sbuffer.scala 134:17]
  wire  _GEN_4024 = line_mask_clean_valid_1 ? _GEN_3000 : _GEN_1976; // @[Sbuffer.scala 134:17]
  wire  _GEN_4025 = line_mask_clean_valid_1 ? _GEN_3001 : _GEN_1977; // @[Sbuffer.scala 134:17]
  wire  _GEN_4026 = line_mask_clean_valid_1 ? _GEN_3002 : _GEN_1978; // @[Sbuffer.scala 134:17]
  wire  _GEN_4027 = line_mask_clean_valid_1 ? _GEN_3003 : _GEN_1979; // @[Sbuffer.scala 134:17]
  wire  _GEN_4028 = line_mask_clean_valid_1 ? _GEN_3004 : _GEN_1980; // @[Sbuffer.scala 134:17]
  wire  _GEN_4029 = line_mask_clean_valid_1 ? _GEN_3005 : _GEN_1981; // @[Sbuffer.scala 134:17]
  wire  _GEN_4030 = line_mask_clean_valid_1 ? _GEN_3006 : _GEN_1982; // @[Sbuffer.scala 134:17]
  wire  _GEN_4031 = line_mask_clean_valid_1 ? _GEN_3007 : _GEN_1983; // @[Sbuffer.scala 134:17]
  wire  _GEN_4032 = line_mask_clean_valid_1 ? _GEN_3008 : _GEN_1984; // @[Sbuffer.scala 134:17]
  wire  _GEN_4033 = line_mask_clean_valid_1 ? _GEN_3009 : _GEN_1985; // @[Sbuffer.scala 134:17]
  wire  _GEN_4034 = line_mask_clean_valid_1 ? _GEN_3010 : _GEN_1986; // @[Sbuffer.scala 134:17]
  wire  _GEN_4035 = line_mask_clean_valid_1 ? _GEN_3011 : _GEN_1987; // @[Sbuffer.scala 134:17]
  wire  _GEN_4036 = line_mask_clean_valid_1 ? _GEN_3012 : _GEN_1988; // @[Sbuffer.scala 134:17]
  wire  _GEN_4037 = line_mask_clean_valid_1 ? _GEN_3013 : _GEN_1989; // @[Sbuffer.scala 134:17]
  wire  _GEN_4038 = line_mask_clean_valid_1 ? _GEN_3014 : _GEN_1990; // @[Sbuffer.scala 134:17]
  wire  _GEN_4039 = line_mask_clean_valid_1 ? _GEN_3015 : _GEN_1991; // @[Sbuffer.scala 134:17]
  wire  _GEN_4040 = line_mask_clean_valid_1 ? _GEN_3016 : _GEN_1992; // @[Sbuffer.scala 134:17]
  wire  _GEN_4041 = line_mask_clean_valid_1 ? _GEN_3017 : _GEN_1993; // @[Sbuffer.scala 134:17]
  wire  _GEN_4042 = line_mask_clean_valid_1 ? _GEN_3018 : _GEN_1994; // @[Sbuffer.scala 134:17]
  wire  _GEN_4043 = line_mask_clean_valid_1 ? _GEN_3019 : _GEN_1995; // @[Sbuffer.scala 134:17]
  wire  _GEN_4044 = line_mask_clean_valid_1 ? _GEN_3020 : _GEN_1996; // @[Sbuffer.scala 134:17]
  wire  _GEN_4045 = line_mask_clean_valid_1 ? _GEN_3021 : _GEN_1997; // @[Sbuffer.scala 134:17]
  wire  _GEN_4046 = line_mask_clean_valid_1 ? _GEN_3022 : _GEN_1998; // @[Sbuffer.scala 134:17]
  wire  _GEN_4047 = line_mask_clean_valid_1 ? _GEN_3023 : _GEN_1999; // @[Sbuffer.scala 134:17]
  wire  _GEN_4048 = line_mask_clean_valid_1 ? _GEN_3024 : _GEN_2000; // @[Sbuffer.scala 134:17]
  wire  _GEN_4049 = line_mask_clean_valid_1 ? _GEN_3025 : _GEN_2001; // @[Sbuffer.scala 134:17]
  wire  _GEN_4050 = line_mask_clean_valid_1 ? _GEN_3026 : _GEN_2002; // @[Sbuffer.scala 134:17]
  wire  _GEN_4051 = line_mask_clean_valid_1 ? _GEN_3027 : _GEN_2003; // @[Sbuffer.scala 134:17]
  wire  _GEN_4052 = line_mask_clean_valid_1 ? _GEN_3028 : _GEN_2004; // @[Sbuffer.scala 134:17]
  wire  _GEN_4053 = line_mask_clean_valid_1 ? _GEN_3029 : _GEN_2005; // @[Sbuffer.scala 134:17]
  wire  _GEN_4054 = line_mask_clean_valid_1 ? _GEN_3030 : _GEN_2006; // @[Sbuffer.scala 134:17]
  wire  _GEN_4055 = line_mask_clean_valid_1 ? _GEN_3031 : _GEN_2007; // @[Sbuffer.scala 134:17]
  wire  _GEN_4056 = line_mask_clean_valid_1 ? _GEN_3032 : _GEN_2008; // @[Sbuffer.scala 134:17]
  wire  _GEN_4057 = line_mask_clean_valid_1 ? _GEN_3033 : _GEN_2009; // @[Sbuffer.scala 134:17]
  wire  _GEN_4058 = line_mask_clean_valid_1 ? _GEN_3034 : _GEN_2010; // @[Sbuffer.scala 134:17]
  wire  _GEN_4059 = line_mask_clean_valid_1 ? _GEN_3035 : _GEN_2011; // @[Sbuffer.scala 134:17]
  wire  _GEN_4060 = line_mask_clean_valid_1 ? _GEN_3036 : _GEN_2012; // @[Sbuffer.scala 134:17]
  wire  _GEN_4061 = line_mask_clean_valid_1 ? _GEN_3037 : _GEN_2013; // @[Sbuffer.scala 134:17]
  wire  _GEN_4062 = line_mask_clean_valid_1 ? _GEN_3038 : _GEN_2014; // @[Sbuffer.scala 134:17]
  wire  _GEN_4063 = line_mask_clean_valid_1 ? _GEN_3039 : _GEN_2015; // @[Sbuffer.scala 134:17]
  wire  _GEN_4064 = line_mask_clean_valid_1 ? _GEN_3040 : _GEN_2016; // @[Sbuffer.scala 134:17]
  wire  _GEN_4065 = line_mask_clean_valid_1 ? _GEN_3041 : _GEN_2017; // @[Sbuffer.scala 134:17]
  wire  _GEN_4066 = line_mask_clean_valid_1 ? _GEN_3042 : _GEN_2018; // @[Sbuffer.scala 134:17]
  wire  _GEN_4067 = line_mask_clean_valid_1 ? _GEN_3043 : _GEN_2019; // @[Sbuffer.scala 134:17]
  wire  _GEN_4068 = line_mask_clean_valid_1 ? _GEN_3044 : _GEN_2020; // @[Sbuffer.scala 134:17]
  wire  _GEN_4069 = line_mask_clean_valid_1 ? _GEN_3045 : _GEN_2021; // @[Sbuffer.scala 134:17]
  wire  _GEN_4070 = line_mask_clean_valid_1 ? _GEN_3046 : _GEN_2022; // @[Sbuffer.scala 134:17]
  wire  _GEN_4071 = line_mask_clean_valid_1 ? _GEN_3047 : _GEN_2023; // @[Sbuffer.scala 134:17]
  wire  _GEN_4072 = line_mask_clean_valid_1 ? _GEN_3048 : _GEN_2024; // @[Sbuffer.scala 134:17]
  wire  _GEN_4073 = line_mask_clean_valid_1 ? _GEN_3049 : _GEN_2025; // @[Sbuffer.scala 134:17]
  wire  _GEN_4074 = line_mask_clean_valid_1 ? _GEN_3050 : _GEN_2026; // @[Sbuffer.scala 134:17]
  wire  _GEN_4075 = line_mask_clean_valid_1 ? _GEN_3051 : _GEN_2027; // @[Sbuffer.scala 134:17]
  wire  _GEN_4076 = line_mask_clean_valid_1 ? _GEN_3052 : _GEN_2028; // @[Sbuffer.scala 134:17]
  wire  _GEN_4077 = line_mask_clean_valid_1 ? _GEN_3053 : _GEN_2029; // @[Sbuffer.scala 134:17]
  wire  _GEN_4078 = line_mask_clean_valid_1 ? _GEN_3054 : _GEN_2030; // @[Sbuffer.scala 134:17]
  wire  _GEN_4079 = line_mask_clean_valid_1 ? _GEN_3055 : _GEN_2031; // @[Sbuffer.scala 134:17]
  wire  _GEN_4080 = line_mask_clean_valid_1 ? _GEN_3056 : _GEN_2032; // @[Sbuffer.scala 134:17]
  wire  _GEN_4081 = line_mask_clean_valid_1 ? _GEN_3057 : _GEN_2033; // @[Sbuffer.scala 134:17]
  wire  _GEN_4082 = line_mask_clean_valid_1 ? _GEN_3058 : _GEN_2034; // @[Sbuffer.scala 134:17]
  wire  _GEN_4083 = line_mask_clean_valid_1 ? _GEN_3059 : _GEN_2035; // @[Sbuffer.scala 134:17]
  wire  _GEN_4084 = line_mask_clean_valid_1 ? _GEN_3060 : _GEN_2036; // @[Sbuffer.scala 134:17]
  wire  _GEN_4085 = line_mask_clean_valid_1 ? _GEN_3061 : _GEN_2037; // @[Sbuffer.scala 134:17]
  wire  _GEN_4086 = line_mask_clean_valid_1 ? _GEN_3062 : _GEN_2038; // @[Sbuffer.scala 134:17]
  wire  _GEN_4087 = line_mask_clean_valid_1 ? _GEN_3063 : _GEN_2039; // @[Sbuffer.scala 134:17]
  wire  _GEN_4088 = line_mask_clean_valid_1 ? _GEN_3064 : _GEN_2040; // @[Sbuffer.scala 134:17]
  wire  _GEN_4089 = line_mask_clean_valid_1 ? _GEN_3065 : _GEN_2041; // @[Sbuffer.scala 134:17]
  wire  _GEN_4090 = line_mask_clean_valid_1 ? _GEN_3066 : _GEN_2042; // @[Sbuffer.scala 134:17]
  wire  _GEN_4091 = line_mask_clean_valid_1 ? _GEN_3067 : _GEN_2043; // @[Sbuffer.scala 134:17]
  wire  _GEN_4092 = line_mask_clean_valid_1 ? _GEN_3068 : _GEN_2044; // @[Sbuffer.scala 134:17]
  wire  _GEN_4093 = line_mask_clean_valid_1 ? _GEN_3069 : _GEN_2045; // @[Sbuffer.scala 134:17]
  wire  _GEN_4094 = line_mask_clean_valid_1 ? _GEN_3070 : _GEN_2046; // @[Sbuffer.scala 134:17]
  wire  _GEN_4095 = line_mask_clean_valid_1 ? _GEN_3071 : _GEN_2047; // @[Sbuffer.scala 134:17]
  reg  w_valid_s1_0; // @[Sbuffer.scala 146:40]
  reg  w_valid_s1_1; // @[Sbuffer.scala 146:40]
  reg [63:0] w_data_s1_0; // @[Sbuffer.scala 147:39]
  reg [63:0] w_data_s1_1; // @[Sbuffer.scala 147:39]
  reg  w_wline_s1_0; // @[Sbuffer.scala 148:40]
  reg  w_wline_s1_1; // @[Sbuffer.scala 148:40]
  reg [7:0] w_mask_s1_0; // @[Sbuffer.scala 149:39]
  reg [7:0] w_mask_s1_1; // @[Sbuffer.scala 149:39]
  wire [7:0] w_addr_s1_hi = io_writeReq_0_bits_wvec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_addr_s1_lo = io_writeReq_0_bits_wvec[7:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T = |w_addr_s1_hi; // @[OneHot.scala 32:14]
  wire [7:0] _w_addr_s1_T_1 = w_addr_s1_hi | w_addr_s1_lo; // @[OneHot.scala 32:28]
  wire [3:0] w_addr_s1_hi_1 = _w_addr_s1_T_1[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_addr_s1_lo_1 = _w_addr_s1_T_1[3:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T_2 = |w_addr_s1_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _w_addr_s1_T_3 = w_addr_s1_hi_1 | w_addr_s1_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] w_addr_s1_hi_2 = _w_addr_s1_T_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_addr_s1_lo_2 = _w_addr_s1_T_3[1:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T_4 = |w_addr_s1_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _w_addr_s1_T_5 = w_addr_s1_hi_2 | w_addr_s1_lo_2; // @[OneHot.scala 32:28]
  wire [2:0] _w_addr_s1_T_8 = {_w_addr_s1_T_2,_w_addr_s1_T_4,_w_addr_s1_T_5[1]}; // @[Cat.scala 33:92]
  reg [3:0] w_addr_s1_0; // @[Sbuffer.scala 150:39]
  wire [7:0] w_addr_s1_hi_3 = io_writeReq_1_bits_wvec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_addr_s1_lo_3 = io_writeReq_1_bits_wvec[7:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T_10 = |w_addr_s1_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _w_addr_s1_T_11 = w_addr_s1_hi_3 | w_addr_s1_lo_3; // @[OneHot.scala 32:28]
  wire [3:0] w_addr_s1_hi_4 = _w_addr_s1_T_11[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_addr_s1_lo_4 = _w_addr_s1_T_11[3:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T_12 = |w_addr_s1_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _w_addr_s1_T_13 = w_addr_s1_hi_4 | w_addr_s1_lo_4; // @[OneHot.scala 32:28]
  wire [1:0] w_addr_s1_hi_5 = _w_addr_s1_T_13[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_addr_s1_lo_5 = _w_addr_s1_T_13[1:0]; // @[OneHot.scala 31:18]
  wire  _w_addr_s1_T_14 = |w_addr_s1_hi_5; // @[OneHot.scala 32:14]
  wire [1:0] _w_addr_s1_T_15 = w_addr_s1_hi_5 | w_addr_s1_lo_5; // @[OneHot.scala 32:28]
  wire [2:0] _w_addr_s1_T_18 = {_w_addr_s1_T_12,_w_addr_s1_T_14,_w_addr_s1_T_15[1]}; // @[Cat.scala 33:92]
  reg [3:0] w_addr_s1_1; // @[Sbuffer.scala 150:39]
  reg [2:0] w_word_offset_s1_0; // @[Sbuffer.scala 151:46]
  reg [2:0] w_word_offset_s1_1; // @[Sbuffer.scala 151:46]
  wire  _wen_T_3 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen = w_valid_s1_0 & _wen_T_3; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4096 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4097 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4098 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4099 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4100 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4101 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4102 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4103 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4104 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4105 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4106 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4107 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4108 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4109 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4110 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4111 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_0_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4112 = 4'h0 == w_addr_s1_0 | _GEN_3072; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4113 = 4'h1 == w_addr_s1_0 | _GEN_3073; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4114 = 4'h2 == w_addr_s1_0 | _GEN_3074; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4115 = 4'h3 == w_addr_s1_0 | _GEN_3075; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4116 = 4'h4 == w_addr_s1_0 | _GEN_3076; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4117 = 4'h5 == w_addr_s1_0 | _GEN_3077; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4118 = 4'h6 == w_addr_s1_0 | _GEN_3078; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4119 = 4'h7 == w_addr_s1_0 | _GEN_3079; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4120 = 4'h8 == w_addr_s1_0 | _GEN_3080; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4121 = 4'h9 == w_addr_s1_0 | _GEN_3081; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4122 = 4'ha == w_addr_s1_0 | _GEN_3082; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4123 = 4'hb == w_addr_s1_0 | _GEN_3083; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4124 = 4'hc == w_addr_s1_0 | _GEN_3084; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4125 = 4'hd == w_addr_s1_0 | _GEN_3085; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4126 = 4'he == w_addr_s1_0 | _GEN_3086; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4127 = 4'hf == w_addr_s1_0 | _GEN_3087; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4128 = wen ? _GEN_4096 : data_0_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4129 = wen ? _GEN_4097 : data_1_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4130 = wen ? _GEN_4098 : data_2_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4131 = wen ? _GEN_4099 : data_3_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4132 = wen ? _GEN_4100 : data_4_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4133 = wen ? _GEN_4101 : data_5_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4134 = wen ? _GEN_4102 : data_6_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4135 = wen ? _GEN_4103 : data_7_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4136 = wen ? _GEN_4104 : data_8_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4137 = wen ? _GEN_4105 : data_9_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4138 = wen ? _GEN_4106 : data_10_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4139 = wen ? _GEN_4107 : data_11_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4140 = wen ? _GEN_4108 : data_12_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4141 = wen ? _GEN_4109 : data_13_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4142 = wen ? _GEN_4110 : data_14_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4143 = wen ? _GEN_4111 : data_15_0_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4144 = wen ? _GEN_4112 : _GEN_3072; // @[Sbuffer.scala 160:18]
  wire  _GEN_4145 = wen ? _GEN_4113 : _GEN_3073; // @[Sbuffer.scala 160:18]
  wire  _GEN_4146 = wen ? _GEN_4114 : _GEN_3074; // @[Sbuffer.scala 160:18]
  wire  _GEN_4147 = wen ? _GEN_4115 : _GEN_3075; // @[Sbuffer.scala 160:18]
  wire  _GEN_4148 = wen ? _GEN_4116 : _GEN_3076; // @[Sbuffer.scala 160:18]
  wire  _GEN_4149 = wen ? _GEN_4117 : _GEN_3077; // @[Sbuffer.scala 160:18]
  wire  _GEN_4150 = wen ? _GEN_4118 : _GEN_3078; // @[Sbuffer.scala 160:18]
  wire  _GEN_4151 = wen ? _GEN_4119 : _GEN_3079; // @[Sbuffer.scala 160:18]
  wire  _GEN_4152 = wen ? _GEN_4120 : _GEN_3080; // @[Sbuffer.scala 160:18]
  wire  _GEN_4153 = wen ? _GEN_4121 : _GEN_3081; // @[Sbuffer.scala 160:18]
  wire  _GEN_4154 = wen ? _GEN_4122 : _GEN_3082; // @[Sbuffer.scala 160:18]
  wire  _GEN_4155 = wen ? _GEN_4123 : _GEN_3083; // @[Sbuffer.scala 160:18]
  wire  _GEN_4156 = wen ? _GEN_4124 : _GEN_3084; // @[Sbuffer.scala 160:18]
  wire  _GEN_4157 = wen ? _GEN_4125 : _GEN_3085; // @[Sbuffer.scala 160:18]
  wire  _GEN_4158 = wen ? _GEN_4126 : _GEN_3086; // @[Sbuffer.scala 160:18]
  wire  _GEN_4159 = wen ? _GEN_4127 : _GEN_3087; // @[Sbuffer.scala 160:18]
  wire  _wen_T_7 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_1 = w_valid_s1_0 & _wen_T_7; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4160 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4161 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4162 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4163 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4164 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4165 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4166 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4167 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4168 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4169 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4170 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4171 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4172 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4173 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4174 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4175 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_0_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4176 = 4'h0 == w_addr_s1_0 | _GEN_3088; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4177 = 4'h1 == w_addr_s1_0 | _GEN_3089; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4178 = 4'h2 == w_addr_s1_0 | _GEN_3090; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4179 = 4'h3 == w_addr_s1_0 | _GEN_3091; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4180 = 4'h4 == w_addr_s1_0 | _GEN_3092; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4181 = 4'h5 == w_addr_s1_0 | _GEN_3093; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4182 = 4'h6 == w_addr_s1_0 | _GEN_3094; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4183 = 4'h7 == w_addr_s1_0 | _GEN_3095; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4184 = 4'h8 == w_addr_s1_0 | _GEN_3096; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4185 = 4'h9 == w_addr_s1_0 | _GEN_3097; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4186 = 4'ha == w_addr_s1_0 | _GEN_3098; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4187 = 4'hb == w_addr_s1_0 | _GEN_3099; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4188 = 4'hc == w_addr_s1_0 | _GEN_3100; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4189 = 4'hd == w_addr_s1_0 | _GEN_3101; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4190 = 4'he == w_addr_s1_0 | _GEN_3102; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4191 = 4'hf == w_addr_s1_0 | _GEN_3103; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4192 = wen_1 ? _GEN_4160 : data_0_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4193 = wen_1 ? _GEN_4161 : data_1_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4194 = wen_1 ? _GEN_4162 : data_2_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4195 = wen_1 ? _GEN_4163 : data_3_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4196 = wen_1 ? _GEN_4164 : data_4_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4197 = wen_1 ? _GEN_4165 : data_5_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4198 = wen_1 ? _GEN_4166 : data_6_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4199 = wen_1 ? _GEN_4167 : data_7_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4200 = wen_1 ? _GEN_4168 : data_8_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4201 = wen_1 ? _GEN_4169 : data_9_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4202 = wen_1 ? _GEN_4170 : data_10_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4203 = wen_1 ? _GEN_4171 : data_11_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4204 = wen_1 ? _GEN_4172 : data_12_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4205 = wen_1 ? _GEN_4173 : data_13_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4206 = wen_1 ? _GEN_4174 : data_14_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4207 = wen_1 ? _GEN_4175 : data_15_0_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4208 = wen_1 ? _GEN_4176 : _GEN_3088; // @[Sbuffer.scala 160:18]
  wire  _GEN_4209 = wen_1 ? _GEN_4177 : _GEN_3089; // @[Sbuffer.scala 160:18]
  wire  _GEN_4210 = wen_1 ? _GEN_4178 : _GEN_3090; // @[Sbuffer.scala 160:18]
  wire  _GEN_4211 = wen_1 ? _GEN_4179 : _GEN_3091; // @[Sbuffer.scala 160:18]
  wire  _GEN_4212 = wen_1 ? _GEN_4180 : _GEN_3092; // @[Sbuffer.scala 160:18]
  wire  _GEN_4213 = wen_1 ? _GEN_4181 : _GEN_3093; // @[Sbuffer.scala 160:18]
  wire  _GEN_4214 = wen_1 ? _GEN_4182 : _GEN_3094; // @[Sbuffer.scala 160:18]
  wire  _GEN_4215 = wen_1 ? _GEN_4183 : _GEN_3095; // @[Sbuffer.scala 160:18]
  wire  _GEN_4216 = wen_1 ? _GEN_4184 : _GEN_3096; // @[Sbuffer.scala 160:18]
  wire  _GEN_4217 = wen_1 ? _GEN_4185 : _GEN_3097; // @[Sbuffer.scala 160:18]
  wire  _GEN_4218 = wen_1 ? _GEN_4186 : _GEN_3098; // @[Sbuffer.scala 160:18]
  wire  _GEN_4219 = wen_1 ? _GEN_4187 : _GEN_3099; // @[Sbuffer.scala 160:18]
  wire  _GEN_4220 = wen_1 ? _GEN_4188 : _GEN_3100; // @[Sbuffer.scala 160:18]
  wire  _GEN_4221 = wen_1 ? _GEN_4189 : _GEN_3101; // @[Sbuffer.scala 160:18]
  wire  _GEN_4222 = wen_1 ? _GEN_4190 : _GEN_3102; // @[Sbuffer.scala 160:18]
  wire  _GEN_4223 = wen_1 ? _GEN_4191 : _GEN_3103; // @[Sbuffer.scala 160:18]
  wire  _wen_T_11 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_2 = w_valid_s1_0 & _wen_T_11; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4224 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4225 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4226 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4227 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4228 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4229 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4230 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4231 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4232 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4233 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4234 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4235 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4236 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4237 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4238 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4239 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_0_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4240 = 4'h0 == w_addr_s1_0 | _GEN_3104; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4241 = 4'h1 == w_addr_s1_0 | _GEN_3105; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4242 = 4'h2 == w_addr_s1_0 | _GEN_3106; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4243 = 4'h3 == w_addr_s1_0 | _GEN_3107; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4244 = 4'h4 == w_addr_s1_0 | _GEN_3108; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4245 = 4'h5 == w_addr_s1_0 | _GEN_3109; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4246 = 4'h6 == w_addr_s1_0 | _GEN_3110; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4247 = 4'h7 == w_addr_s1_0 | _GEN_3111; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4248 = 4'h8 == w_addr_s1_0 | _GEN_3112; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4249 = 4'h9 == w_addr_s1_0 | _GEN_3113; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4250 = 4'ha == w_addr_s1_0 | _GEN_3114; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4251 = 4'hb == w_addr_s1_0 | _GEN_3115; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4252 = 4'hc == w_addr_s1_0 | _GEN_3116; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4253 = 4'hd == w_addr_s1_0 | _GEN_3117; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4254 = 4'he == w_addr_s1_0 | _GEN_3118; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4255 = 4'hf == w_addr_s1_0 | _GEN_3119; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4256 = wen_2 ? _GEN_4224 : data_0_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4257 = wen_2 ? _GEN_4225 : data_1_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4258 = wen_2 ? _GEN_4226 : data_2_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4259 = wen_2 ? _GEN_4227 : data_3_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4260 = wen_2 ? _GEN_4228 : data_4_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4261 = wen_2 ? _GEN_4229 : data_5_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4262 = wen_2 ? _GEN_4230 : data_6_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4263 = wen_2 ? _GEN_4231 : data_7_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4264 = wen_2 ? _GEN_4232 : data_8_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4265 = wen_2 ? _GEN_4233 : data_9_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4266 = wen_2 ? _GEN_4234 : data_10_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4267 = wen_2 ? _GEN_4235 : data_11_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4268 = wen_2 ? _GEN_4236 : data_12_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4269 = wen_2 ? _GEN_4237 : data_13_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4270 = wen_2 ? _GEN_4238 : data_14_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4271 = wen_2 ? _GEN_4239 : data_15_0_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4272 = wen_2 ? _GEN_4240 : _GEN_3104; // @[Sbuffer.scala 160:18]
  wire  _GEN_4273 = wen_2 ? _GEN_4241 : _GEN_3105; // @[Sbuffer.scala 160:18]
  wire  _GEN_4274 = wen_2 ? _GEN_4242 : _GEN_3106; // @[Sbuffer.scala 160:18]
  wire  _GEN_4275 = wen_2 ? _GEN_4243 : _GEN_3107; // @[Sbuffer.scala 160:18]
  wire  _GEN_4276 = wen_2 ? _GEN_4244 : _GEN_3108; // @[Sbuffer.scala 160:18]
  wire  _GEN_4277 = wen_2 ? _GEN_4245 : _GEN_3109; // @[Sbuffer.scala 160:18]
  wire  _GEN_4278 = wen_2 ? _GEN_4246 : _GEN_3110; // @[Sbuffer.scala 160:18]
  wire  _GEN_4279 = wen_2 ? _GEN_4247 : _GEN_3111; // @[Sbuffer.scala 160:18]
  wire  _GEN_4280 = wen_2 ? _GEN_4248 : _GEN_3112; // @[Sbuffer.scala 160:18]
  wire  _GEN_4281 = wen_2 ? _GEN_4249 : _GEN_3113; // @[Sbuffer.scala 160:18]
  wire  _GEN_4282 = wen_2 ? _GEN_4250 : _GEN_3114; // @[Sbuffer.scala 160:18]
  wire  _GEN_4283 = wen_2 ? _GEN_4251 : _GEN_3115; // @[Sbuffer.scala 160:18]
  wire  _GEN_4284 = wen_2 ? _GEN_4252 : _GEN_3116; // @[Sbuffer.scala 160:18]
  wire  _GEN_4285 = wen_2 ? _GEN_4253 : _GEN_3117; // @[Sbuffer.scala 160:18]
  wire  _GEN_4286 = wen_2 ? _GEN_4254 : _GEN_3118; // @[Sbuffer.scala 160:18]
  wire  _GEN_4287 = wen_2 ? _GEN_4255 : _GEN_3119; // @[Sbuffer.scala 160:18]
  wire  _wen_T_15 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_3 = w_valid_s1_0 & _wen_T_15; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4288 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4289 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4290 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4291 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4292 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4293 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4294 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4295 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4296 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4297 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4298 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4299 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4300 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4301 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4302 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4303 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_0_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4304 = 4'h0 == w_addr_s1_0 | _GEN_3120; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4305 = 4'h1 == w_addr_s1_0 | _GEN_3121; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4306 = 4'h2 == w_addr_s1_0 | _GEN_3122; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4307 = 4'h3 == w_addr_s1_0 | _GEN_3123; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4308 = 4'h4 == w_addr_s1_0 | _GEN_3124; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4309 = 4'h5 == w_addr_s1_0 | _GEN_3125; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4310 = 4'h6 == w_addr_s1_0 | _GEN_3126; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4311 = 4'h7 == w_addr_s1_0 | _GEN_3127; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4312 = 4'h8 == w_addr_s1_0 | _GEN_3128; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4313 = 4'h9 == w_addr_s1_0 | _GEN_3129; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4314 = 4'ha == w_addr_s1_0 | _GEN_3130; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4315 = 4'hb == w_addr_s1_0 | _GEN_3131; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4316 = 4'hc == w_addr_s1_0 | _GEN_3132; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4317 = 4'hd == w_addr_s1_0 | _GEN_3133; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4318 = 4'he == w_addr_s1_0 | _GEN_3134; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4319 = 4'hf == w_addr_s1_0 | _GEN_3135; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4320 = wen_3 ? _GEN_4288 : data_0_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4321 = wen_3 ? _GEN_4289 : data_1_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4322 = wen_3 ? _GEN_4290 : data_2_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4323 = wen_3 ? _GEN_4291 : data_3_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4324 = wen_3 ? _GEN_4292 : data_4_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4325 = wen_3 ? _GEN_4293 : data_5_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4326 = wen_3 ? _GEN_4294 : data_6_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4327 = wen_3 ? _GEN_4295 : data_7_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4328 = wen_3 ? _GEN_4296 : data_8_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4329 = wen_3 ? _GEN_4297 : data_9_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4330 = wen_3 ? _GEN_4298 : data_10_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4331 = wen_3 ? _GEN_4299 : data_11_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4332 = wen_3 ? _GEN_4300 : data_12_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4333 = wen_3 ? _GEN_4301 : data_13_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4334 = wen_3 ? _GEN_4302 : data_14_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4335 = wen_3 ? _GEN_4303 : data_15_0_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4336 = wen_3 ? _GEN_4304 : _GEN_3120; // @[Sbuffer.scala 160:18]
  wire  _GEN_4337 = wen_3 ? _GEN_4305 : _GEN_3121; // @[Sbuffer.scala 160:18]
  wire  _GEN_4338 = wen_3 ? _GEN_4306 : _GEN_3122; // @[Sbuffer.scala 160:18]
  wire  _GEN_4339 = wen_3 ? _GEN_4307 : _GEN_3123; // @[Sbuffer.scala 160:18]
  wire  _GEN_4340 = wen_3 ? _GEN_4308 : _GEN_3124; // @[Sbuffer.scala 160:18]
  wire  _GEN_4341 = wen_3 ? _GEN_4309 : _GEN_3125; // @[Sbuffer.scala 160:18]
  wire  _GEN_4342 = wen_3 ? _GEN_4310 : _GEN_3126; // @[Sbuffer.scala 160:18]
  wire  _GEN_4343 = wen_3 ? _GEN_4311 : _GEN_3127; // @[Sbuffer.scala 160:18]
  wire  _GEN_4344 = wen_3 ? _GEN_4312 : _GEN_3128; // @[Sbuffer.scala 160:18]
  wire  _GEN_4345 = wen_3 ? _GEN_4313 : _GEN_3129; // @[Sbuffer.scala 160:18]
  wire  _GEN_4346 = wen_3 ? _GEN_4314 : _GEN_3130; // @[Sbuffer.scala 160:18]
  wire  _GEN_4347 = wen_3 ? _GEN_4315 : _GEN_3131; // @[Sbuffer.scala 160:18]
  wire  _GEN_4348 = wen_3 ? _GEN_4316 : _GEN_3132; // @[Sbuffer.scala 160:18]
  wire  _GEN_4349 = wen_3 ? _GEN_4317 : _GEN_3133; // @[Sbuffer.scala 160:18]
  wire  _GEN_4350 = wen_3 ? _GEN_4318 : _GEN_3134; // @[Sbuffer.scala 160:18]
  wire  _GEN_4351 = wen_3 ? _GEN_4319 : _GEN_3135; // @[Sbuffer.scala 160:18]
  wire  _wen_T_19 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_4 = w_valid_s1_0 & _wen_T_19; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4352 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4353 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4354 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4355 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4356 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4357 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4358 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4359 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4360 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4361 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4362 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4363 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4364 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4365 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4366 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4367 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_0_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4368 = 4'h0 == w_addr_s1_0 | _GEN_3136; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4369 = 4'h1 == w_addr_s1_0 | _GEN_3137; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4370 = 4'h2 == w_addr_s1_0 | _GEN_3138; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4371 = 4'h3 == w_addr_s1_0 | _GEN_3139; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4372 = 4'h4 == w_addr_s1_0 | _GEN_3140; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4373 = 4'h5 == w_addr_s1_0 | _GEN_3141; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4374 = 4'h6 == w_addr_s1_0 | _GEN_3142; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4375 = 4'h7 == w_addr_s1_0 | _GEN_3143; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4376 = 4'h8 == w_addr_s1_0 | _GEN_3144; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4377 = 4'h9 == w_addr_s1_0 | _GEN_3145; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4378 = 4'ha == w_addr_s1_0 | _GEN_3146; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4379 = 4'hb == w_addr_s1_0 | _GEN_3147; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4380 = 4'hc == w_addr_s1_0 | _GEN_3148; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4381 = 4'hd == w_addr_s1_0 | _GEN_3149; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4382 = 4'he == w_addr_s1_0 | _GEN_3150; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4383 = 4'hf == w_addr_s1_0 | _GEN_3151; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4384 = wen_4 ? _GEN_4352 : data_0_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4385 = wen_4 ? _GEN_4353 : data_1_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4386 = wen_4 ? _GEN_4354 : data_2_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4387 = wen_4 ? _GEN_4355 : data_3_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4388 = wen_4 ? _GEN_4356 : data_4_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4389 = wen_4 ? _GEN_4357 : data_5_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4390 = wen_4 ? _GEN_4358 : data_6_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4391 = wen_4 ? _GEN_4359 : data_7_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4392 = wen_4 ? _GEN_4360 : data_8_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4393 = wen_4 ? _GEN_4361 : data_9_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4394 = wen_4 ? _GEN_4362 : data_10_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4395 = wen_4 ? _GEN_4363 : data_11_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4396 = wen_4 ? _GEN_4364 : data_12_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4397 = wen_4 ? _GEN_4365 : data_13_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4398 = wen_4 ? _GEN_4366 : data_14_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4399 = wen_4 ? _GEN_4367 : data_15_0_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4400 = wen_4 ? _GEN_4368 : _GEN_3136; // @[Sbuffer.scala 160:18]
  wire  _GEN_4401 = wen_4 ? _GEN_4369 : _GEN_3137; // @[Sbuffer.scala 160:18]
  wire  _GEN_4402 = wen_4 ? _GEN_4370 : _GEN_3138; // @[Sbuffer.scala 160:18]
  wire  _GEN_4403 = wen_4 ? _GEN_4371 : _GEN_3139; // @[Sbuffer.scala 160:18]
  wire  _GEN_4404 = wen_4 ? _GEN_4372 : _GEN_3140; // @[Sbuffer.scala 160:18]
  wire  _GEN_4405 = wen_4 ? _GEN_4373 : _GEN_3141; // @[Sbuffer.scala 160:18]
  wire  _GEN_4406 = wen_4 ? _GEN_4374 : _GEN_3142; // @[Sbuffer.scala 160:18]
  wire  _GEN_4407 = wen_4 ? _GEN_4375 : _GEN_3143; // @[Sbuffer.scala 160:18]
  wire  _GEN_4408 = wen_4 ? _GEN_4376 : _GEN_3144; // @[Sbuffer.scala 160:18]
  wire  _GEN_4409 = wen_4 ? _GEN_4377 : _GEN_3145; // @[Sbuffer.scala 160:18]
  wire  _GEN_4410 = wen_4 ? _GEN_4378 : _GEN_3146; // @[Sbuffer.scala 160:18]
  wire  _GEN_4411 = wen_4 ? _GEN_4379 : _GEN_3147; // @[Sbuffer.scala 160:18]
  wire  _GEN_4412 = wen_4 ? _GEN_4380 : _GEN_3148; // @[Sbuffer.scala 160:18]
  wire  _GEN_4413 = wen_4 ? _GEN_4381 : _GEN_3149; // @[Sbuffer.scala 160:18]
  wire  _GEN_4414 = wen_4 ? _GEN_4382 : _GEN_3150; // @[Sbuffer.scala 160:18]
  wire  _GEN_4415 = wen_4 ? _GEN_4383 : _GEN_3151; // @[Sbuffer.scala 160:18]
  wire  _wen_T_23 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_5 = w_valid_s1_0 & _wen_T_23; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4416 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4417 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4418 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4419 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4420 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4421 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4422 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4423 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4424 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4425 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4426 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4427 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4428 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4429 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4430 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4431 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_0_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4432 = 4'h0 == w_addr_s1_0 | _GEN_3152; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4433 = 4'h1 == w_addr_s1_0 | _GEN_3153; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4434 = 4'h2 == w_addr_s1_0 | _GEN_3154; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4435 = 4'h3 == w_addr_s1_0 | _GEN_3155; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4436 = 4'h4 == w_addr_s1_0 | _GEN_3156; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4437 = 4'h5 == w_addr_s1_0 | _GEN_3157; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4438 = 4'h6 == w_addr_s1_0 | _GEN_3158; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4439 = 4'h7 == w_addr_s1_0 | _GEN_3159; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4440 = 4'h8 == w_addr_s1_0 | _GEN_3160; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4441 = 4'h9 == w_addr_s1_0 | _GEN_3161; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4442 = 4'ha == w_addr_s1_0 | _GEN_3162; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4443 = 4'hb == w_addr_s1_0 | _GEN_3163; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4444 = 4'hc == w_addr_s1_0 | _GEN_3164; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4445 = 4'hd == w_addr_s1_0 | _GEN_3165; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4446 = 4'he == w_addr_s1_0 | _GEN_3166; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4447 = 4'hf == w_addr_s1_0 | _GEN_3167; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4448 = wen_5 ? _GEN_4416 : data_0_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4449 = wen_5 ? _GEN_4417 : data_1_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4450 = wen_5 ? _GEN_4418 : data_2_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4451 = wen_5 ? _GEN_4419 : data_3_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4452 = wen_5 ? _GEN_4420 : data_4_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4453 = wen_5 ? _GEN_4421 : data_5_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4454 = wen_5 ? _GEN_4422 : data_6_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4455 = wen_5 ? _GEN_4423 : data_7_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4456 = wen_5 ? _GEN_4424 : data_8_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4457 = wen_5 ? _GEN_4425 : data_9_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4458 = wen_5 ? _GEN_4426 : data_10_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4459 = wen_5 ? _GEN_4427 : data_11_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4460 = wen_5 ? _GEN_4428 : data_12_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4461 = wen_5 ? _GEN_4429 : data_13_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4462 = wen_5 ? _GEN_4430 : data_14_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4463 = wen_5 ? _GEN_4431 : data_15_0_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4464 = wen_5 ? _GEN_4432 : _GEN_3152; // @[Sbuffer.scala 160:18]
  wire  _GEN_4465 = wen_5 ? _GEN_4433 : _GEN_3153; // @[Sbuffer.scala 160:18]
  wire  _GEN_4466 = wen_5 ? _GEN_4434 : _GEN_3154; // @[Sbuffer.scala 160:18]
  wire  _GEN_4467 = wen_5 ? _GEN_4435 : _GEN_3155; // @[Sbuffer.scala 160:18]
  wire  _GEN_4468 = wen_5 ? _GEN_4436 : _GEN_3156; // @[Sbuffer.scala 160:18]
  wire  _GEN_4469 = wen_5 ? _GEN_4437 : _GEN_3157; // @[Sbuffer.scala 160:18]
  wire  _GEN_4470 = wen_5 ? _GEN_4438 : _GEN_3158; // @[Sbuffer.scala 160:18]
  wire  _GEN_4471 = wen_5 ? _GEN_4439 : _GEN_3159; // @[Sbuffer.scala 160:18]
  wire  _GEN_4472 = wen_5 ? _GEN_4440 : _GEN_3160; // @[Sbuffer.scala 160:18]
  wire  _GEN_4473 = wen_5 ? _GEN_4441 : _GEN_3161; // @[Sbuffer.scala 160:18]
  wire  _GEN_4474 = wen_5 ? _GEN_4442 : _GEN_3162; // @[Sbuffer.scala 160:18]
  wire  _GEN_4475 = wen_5 ? _GEN_4443 : _GEN_3163; // @[Sbuffer.scala 160:18]
  wire  _GEN_4476 = wen_5 ? _GEN_4444 : _GEN_3164; // @[Sbuffer.scala 160:18]
  wire  _GEN_4477 = wen_5 ? _GEN_4445 : _GEN_3165; // @[Sbuffer.scala 160:18]
  wire  _GEN_4478 = wen_5 ? _GEN_4446 : _GEN_3166; // @[Sbuffer.scala 160:18]
  wire  _GEN_4479 = wen_5 ? _GEN_4447 : _GEN_3167; // @[Sbuffer.scala 160:18]
  wire  _wen_T_27 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_6 = w_valid_s1_0 & _wen_T_27; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4480 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4481 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4482 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4483 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4484 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4485 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4486 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4487 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4488 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4489 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4490 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4491 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4492 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4493 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4494 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4495 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_0_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4496 = 4'h0 == w_addr_s1_0 | _GEN_3168; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4497 = 4'h1 == w_addr_s1_0 | _GEN_3169; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4498 = 4'h2 == w_addr_s1_0 | _GEN_3170; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4499 = 4'h3 == w_addr_s1_0 | _GEN_3171; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4500 = 4'h4 == w_addr_s1_0 | _GEN_3172; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4501 = 4'h5 == w_addr_s1_0 | _GEN_3173; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4502 = 4'h6 == w_addr_s1_0 | _GEN_3174; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4503 = 4'h7 == w_addr_s1_0 | _GEN_3175; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4504 = 4'h8 == w_addr_s1_0 | _GEN_3176; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4505 = 4'h9 == w_addr_s1_0 | _GEN_3177; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4506 = 4'ha == w_addr_s1_0 | _GEN_3178; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4507 = 4'hb == w_addr_s1_0 | _GEN_3179; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4508 = 4'hc == w_addr_s1_0 | _GEN_3180; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4509 = 4'hd == w_addr_s1_0 | _GEN_3181; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4510 = 4'he == w_addr_s1_0 | _GEN_3182; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4511 = 4'hf == w_addr_s1_0 | _GEN_3183; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4512 = wen_6 ? _GEN_4480 : data_0_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4513 = wen_6 ? _GEN_4481 : data_1_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4514 = wen_6 ? _GEN_4482 : data_2_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4515 = wen_6 ? _GEN_4483 : data_3_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4516 = wen_6 ? _GEN_4484 : data_4_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4517 = wen_6 ? _GEN_4485 : data_5_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4518 = wen_6 ? _GEN_4486 : data_6_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4519 = wen_6 ? _GEN_4487 : data_7_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4520 = wen_6 ? _GEN_4488 : data_8_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4521 = wen_6 ? _GEN_4489 : data_9_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4522 = wen_6 ? _GEN_4490 : data_10_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4523 = wen_6 ? _GEN_4491 : data_11_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4524 = wen_6 ? _GEN_4492 : data_12_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4525 = wen_6 ? _GEN_4493 : data_13_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4526 = wen_6 ? _GEN_4494 : data_14_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4527 = wen_6 ? _GEN_4495 : data_15_0_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4528 = wen_6 ? _GEN_4496 : _GEN_3168; // @[Sbuffer.scala 160:18]
  wire  _GEN_4529 = wen_6 ? _GEN_4497 : _GEN_3169; // @[Sbuffer.scala 160:18]
  wire  _GEN_4530 = wen_6 ? _GEN_4498 : _GEN_3170; // @[Sbuffer.scala 160:18]
  wire  _GEN_4531 = wen_6 ? _GEN_4499 : _GEN_3171; // @[Sbuffer.scala 160:18]
  wire  _GEN_4532 = wen_6 ? _GEN_4500 : _GEN_3172; // @[Sbuffer.scala 160:18]
  wire  _GEN_4533 = wen_6 ? _GEN_4501 : _GEN_3173; // @[Sbuffer.scala 160:18]
  wire  _GEN_4534 = wen_6 ? _GEN_4502 : _GEN_3174; // @[Sbuffer.scala 160:18]
  wire  _GEN_4535 = wen_6 ? _GEN_4503 : _GEN_3175; // @[Sbuffer.scala 160:18]
  wire  _GEN_4536 = wen_6 ? _GEN_4504 : _GEN_3176; // @[Sbuffer.scala 160:18]
  wire  _GEN_4537 = wen_6 ? _GEN_4505 : _GEN_3177; // @[Sbuffer.scala 160:18]
  wire  _GEN_4538 = wen_6 ? _GEN_4506 : _GEN_3178; // @[Sbuffer.scala 160:18]
  wire  _GEN_4539 = wen_6 ? _GEN_4507 : _GEN_3179; // @[Sbuffer.scala 160:18]
  wire  _GEN_4540 = wen_6 ? _GEN_4508 : _GEN_3180; // @[Sbuffer.scala 160:18]
  wire  _GEN_4541 = wen_6 ? _GEN_4509 : _GEN_3181; // @[Sbuffer.scala 160:18]
  wire  _GEN_4542 = wen_6 ? _GEN_4510 : _GEN_3182; // @[Sbuffer.scala 160:18]
  wire  _GEN_4543 = wen_6 ? _GEN_4511 : _GEN_3183; // @[Sbuffer.scala 160:18]
  wire  _wen_T_31 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h0 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_7 = w_valid_s1_0 & _wen_T_31; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4544 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4545 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4546 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4547 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4548 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4549 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4550 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4551 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4552 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4553 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4554 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4555 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4556 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4557 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4558 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4559 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_0_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4560 = 4'h0 == w_addr_s1_0 | _GEN_3184; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4561 = 4'h1 == w_addr_s1_0 | _GEN_3185; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4562 = 4'h2 == w_addr_s1_0 | _GEN_3186; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4563 = 4'h3 == w_addr_s1_0 | _GEN_3187; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4564 = 4'h4 == w_addr_s1_0 | _GEN_3188; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4565 = 4'h5 == w_addr_s1_0 | _GEN_3189; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4566 = 4'h6 == w_addr_s1_0 | _GEN_3190; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4567 = 4'h7 == w_addr_s1_0 | _GEN_3191; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4568 = 4'h8 == w_addr_s1_0 | _GEN_3192; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4569 = 4'h9 == w_addr_s1_0 | _GEN_3193; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4570 = 4'ha == w_addr_s1_0 | _GEN_3194; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4571 = 4'hb == w_addr_s1_0 | _GEN_3195; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4572 = 4'hc == w_addr_s1_0 | _GEN_3196; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4573 = 4'hd == w_addr_s1_0 | _GEN_3197; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4574 = 4'he == w_addr_s1_0 | _GEN_3198; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4575 = 4'hf == w_addr_s1_0 | _GEN_3199; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4576 = wen_7 ? _GEN_4544 : data_0_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4577 = wen_7 ? _GEN_4545 : data_1_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4578 = wen_7 ? _GEN_4546 : data_2_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4579 = wen_7 ? _GEN_4547 : data_3_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4580 = wen_7 ? _GEN_4548 : data_4_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4581 = wen_7 ? _GEN_4549 : data_5_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4582 = wen_7 ? _GEN_4550 : data_6_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4583 = wen_7 ? _GEN_4551 : data_7_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4584 = wen_7 ? _GEN_4552 : data_8_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4585 = wen_7 ? _GEN_4553 : data_9_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4586 = wen_7 ? _GEN_4554 : data_10_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4587 = wen_7 ? _GEN_4555 : data_11_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4588 = wen_7 ? _GEN_4556 : data_12_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4589 = wen_7 ? _GEN_4557 : data_13_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4590 = wen_7 ? _GEN_4558 : data_14_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4591 = wen_7 ? _GEN_4559 : data_15_0_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4592 = wen_7 ? _GEN_4560 : _GEN_3184; // @[Sbuffer.scala 160:18]
  wire  _GEN_4593 = wen_7 ? _GEN_4561 : _GEN_3185; // @[Sbuffer.scala 160:18]
  wire  _GEN_4594 = wen_7 ? _GEN_4562 : _GEN_3186; // @[Sbuffer.scala 160:18]
  wire  _GEN_4595 = wen_7 ? _GEN_4563 : _GEN_3187; // @[Sbuffer.scala 160:18]
  wire  _GEN_4596 = wen_7 ? _GEN_4564 : _GEN_3188; // @[Sbuffer.scala 160:18]
  wire  _GEN_4597 = wen_7 ? _GEN_4565 : _GEN_3189; // @[Sbuffer.scala 160:18]
  wire  _GEN_4598 = wen_7 ? _GEN_4566 : _GEN_3190; // @[Sbuffer.scala 160:18]
  wire  _GEN_4599 = wen_7 ? _GEN_4567 : _GEN_3191; // @[Sbuffer.scala 160:18]
  wire  _GEN_4600 = wen_7 ? _GEN_4568 : _GEN_3192; // @[Sbuffer.scala 160:18]
  wire  _GEN_4601 = wen_7 ? _GEN_4569 : _GEN_3193; // @[Sbuffer.scala 160:18]
  wire  _GEN_4602 = wen_7 ? _GEN_4570 : _GEN_3194; // @[Sbuffer.scala 160:18]
  wire  _GEN_4603 = wen_7 ? _GEN_4571 : _GEN_3195; // @[Sbuffer.scala 160:18]
  wire  _GEN_4604 = wen_7 ? _GEN_4572 : _GEN_3196; // @[Sbuffer.scala 160:18]
  wire  _GEN_4605 = wen_7 ? _GEN_4573 : _GEN_3197; // @[Sbuffer.scala 160:18]
  wire  _GEN_4606 = wen_7 ? _GEN_4574 : _GEN_3198; // @[Sbuffer.scala 160:18]
  wire  _GEN_4607 = wen_7 ? _GEN_4575 : _GEN_3199; // @[Sbuffer.scala 160:18]
  wire  _wen_T_35 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_8 = w_valid_s1_0 & _wen_T_35; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4608 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4609 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4610 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4611 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4612 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4613 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4614 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4615 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4616 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4617 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4618 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4619 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4620 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4621 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4622 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4623 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_1_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4624 = 4'h0 == w_addr_s1_0 | _GEN_3200; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4625 = 4'h1 == w_addr_s1_0 | _GEN_3201; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4626 = 4'h2 == w_addr_s1_0 | _GEN_3202; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4627 = 4'h3 == w_addr_s1_0 | _GEN_3203; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4628 = 4'h4 == w_addr_s1_0 | _GEN_3204; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4629 = 4'h5 == w_addr_s1_0 | _GEN_3205; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4630 = 4'h6 == w_addr_s1_0 | _GEN_3206; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4631 = 4'h7 == w_addr_s1_0 | _GEN_3207; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4632 = 4'h8 == w_addr_s1_0 | _GEN_3208; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4633 = 4'h9 == w_addr_s1_0 | _GEN_3209; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4634 = 4'ha == w_addr_s1_0 | _GEN_3210; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4635 = 4'hb == w_addr_s1_0 | _GEN_3211; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4636 = 4'hc == w_addr_s1_0 | _GEN_3212; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4637 = 4'hd == w_addr_s1_0 | _GEN_3213; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4638 = 4'he == w_addr_s1_0 | _GEN_3214; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4639 = 4'hf == w_addr_s1_0 | _GEN_3215; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4640 = wen_8 ? _GEN_4608 : data_0_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4641 = wen_8 ? _GEN_4609 : data_1_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4642 = wen_8 ? _GEN_4610 : data_2_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4643 = wen_8 ? _GEN_4611 : data_3_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4644 = wen_8 ? _GEN_4612 : data_4_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4645 = wen_8 ? _GEN_4613 : data_5_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4646 = wen_8 ? _GEN_4614 : data_6_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4647 = wen_8 ? _GEN_4615 : data_7_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4648 = wen_8 ? _GEN_4616 : data_8_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4649 = wen_8 ? _GEN_4617 : data_9_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4650 = wen_8 ? _GEN_4618 : data_10_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4651 = wen_8 ? _GEN_4619 : data_11_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4652 = wen_8 ? _GEN_4620 : data_12_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4653 = wen_8 ? _GEN_4621 : data_13_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4654 = wen_8 ? _GEN_4622 : data_14_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4655 = wen_8 ? _GEN_4623 : data_15_1_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4656 = wen_8 ? _GEN_4624 : _GEN_3200; // @[Sbuffer.scala 160:18]
  wire  _GEN_4657 = wen_8 ? _GEN_4625 : _GEN_3201; // @[Sbuffer.scala 160:18]
  wire  _GEN_4658 = wen_8 ? _GEN_4626 : _GEN_3202; // @[Sbuffer.scala 160:18]
  wire  _GEN_4659 = wen_8 ? _GEN_4627 : _GEN_3203; // @[Sbuffer.scala 160:18]
  wire  _GEN_4660 = wen_8 ? _GEN_4628 : _GEN_3204; // @[Sbuffer.scala 160:18]
  wire  _GEN_4661 = wen_8 ? _GEN_4629 : _GEN_3205; // @[Sbuffer.scala 160:18]
  wire  _GEN_4662 = wen_8 ? _GEN_4630 : _GEN_3206; // @[Sbuffer.scala 160:18]
  wire  _GEN_4663 = wen_8 ? _GEN_4631 : _GEN_3207; // @[Sbuffer.scala 160:18]
  wire  _GEN_4664 = wen_8 ? _GEN_4632 : _GEN_3208; // @[Sbuffer.scala 160:18]
  wire  _GEN_4665 = wen_8 ? _GEN_4633 : _GEN_3209; // @[Sbuffer.scala 160:18]
  wire  _GEN_4666 = wen_8 ? _GEN_4634 : _GEN_3210; // @[Sbuffer.scala 160:18]
  wire  _GEN_4667 = wen_8 ? _GEN_4635 : _GEN_3211; // @[Sbuffer.scala 160:18]
  wire  _GEN_4668 = wen_8 ? _GEN_4636 : _GEN_3212; // @[Sbuffer.scala 160:18]
  wire  _GEN_4669 = wen_8 ? _GEN_4637 : _GEN_3213; // @[Sbuffer.scala 160:18]
  wire  _GEN_4670 = wen_8 ? _GEN_4638 : _GEN_3214; // @[Sbuffer.scala 160:18]
  wire  _GEN_4671 = wen_8 ? _GEN_4639 : _GEN_3215; // @[Sbuffer.scala 160:18]
  wire  _wen_T_39 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_9 = w_valid_s1_0 & _wen_T_39; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4672 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4673 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4674 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4675 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4676 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4677 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4678 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4679 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4680 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4681 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4682 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4683 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4684 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4685 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4686 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4687 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_1_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4688 = 4'h0 == w_addr_s1_0 | _GEN_3216; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4689 = 4'h1 == w_addr_s1_0 | _GEN_3217; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4690 = 4'h2 == w_addr_s1_0 | _GEN_3218; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4691 = 4'h3 == w_addr_s1_0 | _GEN_3219; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4692 = 4'h4 == w_addr_s1_0 | _GEN_3220; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4693 = 4'h5 == w_addr_s1_0 | _GEN_3221; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4694 = 4'h6 == w_addr_s1_0 | _GEN_3222; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4695 = 4'h7 == w_addr_s1_0 | _GEN_3223; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4696 = 4'h8 == w_addr_s1_0 | _GEN_3224; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4697 = 4'h9 == w_addr_s1_0 | _GEN_3225; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4698 = 4'ha == w_addr_s1_0 | _GEN_3226; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4699 = 4'hb == w_addr_s1_0 | _GEN_3227; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4700 = 4'hc == w_addr_s1_0 | _GEN_3228; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4701 = 4'hd == w_addr_s1_0 | _GEN_3229; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4702 = 4'he == w_addr_s1_0 | _GEN_3230; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4703 = 4'hf == w_addr_s1_0 | _GEN_3231; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4704 = wen_9 ? _GEN_4672 : data_0_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4705 = wen_9 ? _GEN_4673 : data_1_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4706 = wen_9 ? _GEN_4674 : data_2_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4707 = wen_9 ? _GEN_4675 : data_3_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4708 = wen_9 ? _GEN_4676 : data_4_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4709 = wen_9 ? _GEN_4677 : data_5_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4710 = wen_9 ? _GEN_4678 : data_6_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4711 = wen_9 ? _GEN_4679 : data_7_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4712 = wen_9 ? _GEN_4680 : data_8_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4713 = wen_9 ? _GEN_4681 : data_9_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4714 = wen_9 ? _GEN_4682 : data_10_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4715 = wen_9 ? _GEN_4683 : data_11_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4716 = wen_9 ? _GEN_4684 : data_12_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4717 = wen_9 ? _GEN_4685 : data_13_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4718 = wen_9 ? _GEN_4686 : data_14_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4719 = wen_9 ? _GEN_4687 : data_15_1_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4720 = wen_9 ? _GEN_4688 : _GEN_3216; // @[Sbuffer.scala 160:18]
  wire  _GEN_4721 = wen_9 ? _GEN_4689 : _GEN_3217; // @[Sbuffer.scala 160:18]
  wire  _GEN_4722 = wen_9 ? _GEN_4690 : _GEN_3218; // @[Sbuffer.scala 160:18]
  wire  _GEN_4723 = wen_9 ? _GEN_4691 : _GEN_3219; // @[Sbuffer.scala 160:18]
  wire  _GEN_4724 = wen_9 ? _GEN_4692 : _GEN_3220; // @[Sbuffer.scala 160:18]
  wire  _GEN_4725 = wen_9 ? _GEN_4693 : _GEN_3221; // @[Sbuffer.scala 160:18]
  wire  _GEN_4726 = wen_9 ? _GEN_4694 : _GEN_3222; // @[Sbuffer.scala 160:18]
  wire  _GEN_4727 = wen_9 ? _GEN_4695 : _GEN_3223; // @[Sbuffer.scala 160:18]
  wire  _GEN_4728 = wen_9 ? _GEN_4696 : _GEN_3224; // @[Sbuffer.scala 160:18]
  wire  _GEN_4729 = wen_9 ? _GEN_4697 : _GEN_3225; // @[Sbuffer.scala 160:18]
  wire  _GEN_4730 = wen_9 ? _GEN_4698 : _GEN_3226; // @[Sbuffer.scala 160:18]
  wire  _GEN_4731 = wen_9 ? _GEN_4699 : _GEN_3227; // @[Sbuffer.scala 160:18]
  wire  _GEN_4732 = wen_9 ? _GEN_4700 : _GEN_3228; // @[Sbuffer.scala 160:18]
  wire  _GEN_4733 = wen_9 ? _GEN_4701 : _GEN_3229; // @[Sbuffer.scala 160:18]
  wire  _GEN_4734 = wen_9 ? _GEN_4702 : _GEN_3230; // @[Sbuffer.scala 160:18]
  wire  _GEN_4735 = wen_9 ? _GEN_4703 : _GEN_3231; // @[Sbuffer.scala 160:18]
  wire  _wen_T_43 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_10 = w_valid_s1_0 & _wen_T_43; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4736 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4737 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4738 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4739 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4740 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4741 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4742 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4743 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4744 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4745 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4746 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4747 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4748 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4749 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4750 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4751 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_1_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4752 = 4'h0 == w_addr_s1_0 | _GEN_3232; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4753 = 4'h1 == w_addr_s1_0 | _GEN_3233; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4754 = 4'h2 == w_addr_s1_0 | _GEN_3234; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4755 = 4'h3 == w_addr_s1_0 | _GEN_3235; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4756 = 4'h4 == w_addr_s1_0 | _GEN_3236; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4757 = 4'h5 == w_addr_s1_0 | _GEN_3237; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4758 = 4'h6 == w_addr_s1_0 | _GEN_3238; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4759 = 4'h7 == w_addr_s1_0 | _GEN_3239; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4760 = 4'h8 == w_addr_s1_0 | _GEN_3240; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4761 = 4'h9 == w_addr_s1_0 | _GEN_3241; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4762 = 4'ha == w_addr_s1_0 | _GEN_3242; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4763 = 4'hb == w_addr_s1_0 | _GEN_3243; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4764 = 4'hc == w_addr_s1_0 | _GEN_3244; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4765 = 4'hd == w_addr_s1_0 | _GEN_3245; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4766 = 4'he == w_addr_s1_0 | _GEN_3246; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4767 = 4'hf == w_addr_s1_0 | _GEN_3247; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4768 = wen_10 ? _GEN_4736 : data_0_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4769 = wen_10 ? _GEN_4737 : data_1_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4770 = wen_10 ? _GEN_4738 : data_2_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4771 = wen_10 ? _GEN_4739 : data_3_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4772 = wen_10 ? _GEN_4740 : data_4_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4773 = wen_10 ? _GEN_4741 : data_5_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4774 = wen_10 ? _GEN_4742 : data_6_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4775 = wen_10 ? _GEN_4743 : data_7_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4776 = wen_10 ? _GEN_4744 : data_8_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4777 = wen_10 ? _GEN_4745 : data_9_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4778 = wen_10 ? _GEN_4746 : data_10_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4779 = wen_10 ? _GEN_4747 : data_11_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4780 = wen_10 ? _GEN_4748 : data_12_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4781 = wen_10 ? _GEN_4749 : data_13_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4782 = wen_10 ? _GEN_4750 : data_14_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4783 = wen_10 ? _GEN_4751 : data_15_1_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4784 = wen_10 ? _GEN_4752 : _GEN_3232; // @[Sbuffer.scala 160:18]
  wire  _GEN_4785 = wen_10 ? _GEN_4753 : _GEN_3233; // @[Sbuffer.scala 160:18]
  wire  _GEN_4786 = wen_10 ? _GEN_4754 : _GEN_3234; // @[Sbuffer.scala 160:18]
  wire  _GEN_4787 = wen_10 ? _GEN_4755 : _GEN_3235; // @[Sbuffer.scala 160:18]
  wire  _GEN_4788 = wen_10 ? _GEN_4756 : _GEN_3236; // @[Sbuffer.scala 160:18]
  wire  _GEN_4789 = wen_10 ? _GEN_4757 : _GEN_3237; // @[Sbuffer.scala 160:18]
  wire  _GEN_4790 = wen_10 ? _GEN_4758 : _GEN_3238; // @[Sbuffer.scala 160:18]
  wire  _GEN_4791 = wen_10 ? _GEN_4759 : _GEN_3239; // @[Sbuffer.scala 160:18]
  wire  _GEN_4792 = wen_10 ? _GEN_4760 : _GEN_3240; // @[Sbuffer.scala 160:18]
  wire  _GEN_4793 = wen_10 ? _GEN_4761 : _GEN_3241; // @[Sbuffer.scala 160:18]
  wire  _GEN_4794 = wen_10 ? _GEN_4762 : _GEN_3242; // @[Sbuffer.scala 160:18]
  wire  _GEN_4795 = wen_10 ? _GEN_4763 : _GEN_3243; // @[Sbuffer.scala 160:18]
  wire  _GEN_4796 = wen_10 ? _GEN_4764 : _GEN_3244; // @[Sbuffer.scala 160:18]
  wire  _GEN_4797 = wen_10 ? _GEN_4765 : _GEN_3245; // @[Sbuffer.scala 160:18]
  wire  _GEN_4798 = wen_10 ? _GEN_4766 : _GEN_3246; // @[Sbuffer.scala 160:18]
  wire  _GEN_4799 = wen_10 ? _GEN_4767 : _GEN_3247; // @[Sbuffer.scala 160:18]
  wire  _wen_T_47 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_11 = w_valid_s1_0 & _wen_T_47; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4800 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4801 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4802 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4803 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4804 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4805 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4806 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4807 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4808 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4809 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4810 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4811 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4812 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4813 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4814 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4815 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_1_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4816 = 4'h0 == w_addr_s1_0 | _GEN_3248; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4817 = 4'h1 == w_addr_s1_0 | _GEN_3249; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4818 = 4'h2 == w_addr_s1_0 | _GEN_3250; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4819 = 4'h3 == w_addr_s1_0 | _GEN_3251; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4820 = 4'h4 == w_addr_s1_0 | _GEN_3252; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4821 = 4'h5 == w_addr_s1_0 | _GEN_3253; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4822 = 4'h6 == w_addr_s1_0 | _GEN_3254; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4823 = 4'h7 == w_addr_s1_0 | _GEN_3255; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4824 = 4'h8 == w_addr_s1_0 | _GEN_3256; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4825 = 4'h9 == w_addr_s1_0 | _GEN_3257; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4826 = 4'ha == w_addr_s1_0 | _GEN_3258; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4827 = 4'hb == w_addr_s1_0 | _GEN_3259; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4828 = 4'hc == w_addr_s1_0 | _GEN_3260; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4829 = 4'hd == w_addr_s1_0 | _GEN_3261; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4830 = 4'he == w_addr_s1_0 | _GEN_3262; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4831 = 4'hf == w_addr_s1_0 | _GEN_3263; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4832 = wen_11 ? _GEN_4800 : data_0_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4833 = wen_11 ? _GEN_4801 : data_1_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4834 = wen_11 ? _GEN_4802 : data_2_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4835 = wen_11 ? _GEN_4803 : data_3_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4836 = wen_11 ? _GEN_4804 : data_4_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4837 = wen_11 ? _GEN_4805 : data_5_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4838 = wen_11 ? _GEN_4806 : data_6_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4839 = wen_11 ? _GEN_4807 : data_7_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4840 = wen_11 ? _GEN_4808 : data_8_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4841 = wen_11 ? _GEN_4809 : data_9_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4842 = wen_11 ? _GEN_4810 : data_10_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4843 = wen_11 ? _GEN_4811 : data_11_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4844 = wen_11 ? _GEN_4812 : data_12_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4845 = wen_11 ? _GEN_4813 : data_13_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4846 = wen_11 ? _GEN_4814 : data_14_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4847 = wen_11 ? _GEN_4815 : data_15_1_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4848 = wen_11 ? _GEN_4816 : _GEN_3248; // @[Sbuffer.scala 160:18]
  wire  _GEN_4849 = wen_11 ? _GEN_4817 : _GEN_3249; // @[Sbuffer.scala 160:18]
  wire  _GEN_4850 = wen_11 ? _GEN_4818 : _GEN_3250; // @[Sbuffer.scala 160:18]
  wire  _GEN_4851 = wen_11 ? _GEN_4819 : _GEN_3251; // @[Sbuffer.scala 160:18]
  wire  _GEN_4852 = wen_11 ? _GEN_4820 : _GEN_3252; // @[Sbuffer.scala 160:18]
  wire  _GEN_4853 = wen_11 ? _GEN_4821 : _GEN_3253; // @[Sbuffer.scala 160:18]
  wire  _GEN_4854 = wen_11 ? _GEN_4822 : _GEN_3254; // @[Sbuffer.scala 160:18]
  wire  _GEN_4855 = wen_11 ? _GEN_4823 : _GEN_3255; // @[Sbuffer.scala 160:18]
  wire  _GEN_4856 = wen_11 ? _GEN_4824 : _GEN_3256; // @[Sbuffer.scala 160:18]
  wire  _GEN_4857 = wen_11 ? _GEN_4825 : _GEN_3257; // @[Sbuffer.scala 160:18]
  wire  _GEN_4858 = wen_11 ? _GEN_4826 : _GEN_3258; // @[Sbuffer.scala 160:18]
  wire  _GEN_4859 = wen_11 ? _GEN_4827 : _GEN_3259; // @[Sbuffer.scala 160:18]
  wire  _GEN_4860 = wen_11 ? _GEN_4828 : _GEN_3260; // @[Sbuffer.scala 160:18]
  wire  _GEN_4861 = wen_11 ? _GEN_4829 : _GEN_3261; // @[Sbuffer.scala 160:18]
  wire  _GEN_4862 = wen_11 ? _GEN_4830 : _GEN_3262; // @[Sbuffer.scala 160:18]
  wire  _GEN_4863 = wen_11 ? _GEN_4831 : _GEN_3263; // @[Sbuffer.scala 160:18]
  wire  _wen_T_51 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_12 = w_valid_s1_0 & _wen_T_51; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4864 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4865 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4866 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4867 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4868 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4869 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4870 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4871 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4872 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4873 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4874 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4875 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4876 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4877 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4878 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4879 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_1_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4880 = 4'h0 == w_addr_s1_0 | _GEN_3264; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4881 = 4'h1 == w_addr_s1_0 | _GEN_3265; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4882 = 4'h2 == w_addr_s1_0 | _GEN_3266; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4883 = 4'h3 == w_addr_s1_0 | _GEN_3267; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4884 = 4'h4 == w_addr_s1_0 | _GEN_3268; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4885 = 4'h5 == w_addr_s1_0 | _GEN_3269; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4886 = 4'h6 == w_addr_s1_0 | _GEN_3270; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4887 = 4'h7 == w_addr_s1_0 | _GEN_3271; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4888 = 4'h8 == w_addr_s1_0 | _GEN_3272; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4889 = 4'h9 == w_addr_s1_0 | _GEN_3273; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4890 = 4'ha == w_addr_s1_0 | _GEN_3274; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4891 = 4'hb == w_addr_s1_0 | _GEN_3275; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4892 = 4'hc == w_addr_s1_0 | _GEN_3276; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4893 = 4'hd == w_addr_s1_0 | _GEN_3277; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4894 = 4'he == w_addr_s1_0 | _GEN_3278; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4895 = 4'hf == w_addr_s1_0 | _GEN_3279; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4896 = wen_12 ? _GEN_4864 : data_0_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4897 = wen_12 ? _GEN_4865 : data_1_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4898 = wen_12 ? _GEN_4866 : data_2_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4899 = wen_12 ? _GEN_4867 : data_3_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4900 = wen_12 ? _GEN_4868 : data_4_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4901 = wen_12 ? _GEN_4869 : data_5_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4902 = wen_12 ? _GEN_4870 : data_6_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4903 = wen_12 ? _GEN_4871 : data_7_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4904 = wen_12 ? _GEN_4872 : data_8_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4905 = wen_12 ? _GEN_4873 : data_9_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4906 = wen_12 ? _GEN_4874 : data_10_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4907 = wen_12 ? _GEN_4875 : data_11_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4908 = wen_12 ? _GEN_4876 : data_12_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4909 = wen_12 ? _GEN_4877 : data_13_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4910 = wen_12 ? _GEN_4878 : data_14_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4911 = wen_12 ? _GEN_4879 : data_15_1_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4912 = wen_12 ? _GEN_4880 : _GEN_3264; // @[Sbuffer.scala 160:18]
  wire  _GEN_4913 = wen_12 ? _GEN_4881 : _GEN_3265; // @[Sbuffer.scala 160:18]
  wire  _GEN_4914 = wen_12 ? _GEN_4882 : _GEN_3266; // @[Sbuffer.scala 160:18]
  wire  _GEN_4915 = wen_12 ? _GEN_4883 : _GEN_3267; // @[Sbuffer.scala 160:18]
  wire  _GEN_4916 = wen_12 ? _GEN_4884 : _GEN_3268; // @[Sbuffer.scala 160:18]
  wire  _GEN_4917 = wen_12 ? _GEN_4885 : _GEN_3269; // @[Sbuffer.scala 160:18]
  wire  _GEN_4918 = wen_12 ? _GEN_4886 : _GEN_3270; // @[Sbuffer.scala 160:18]
  wire  _GEN_4919 = wen_12 ? _GEN_4887 : _GEN_3271; // @[Sbuffer.scala 160:18]
  wire  _GEN_4920 = wen_12 ? _GEN_4888 : _GEN_3272; // @[Sbuffer.scala 160:18]
  wire  _GEN_4921 = wen_12 ? _GEN_4889 : _GEN_3273; // @[Sbuffer.scala 160:18]
  wire  _GEN_4922 = wen_12 ? _GEN_4890 : _GEN_3274; // @[Sbuffer.scala 160:18]
  wire  _GEN_4923 = wen_12 ? _GEN_4891 : _GEN_3275; // @[Sbuffer.scala 160:18]
  wire  _GEN_4924 = wen_12 ? _GEN_4892 : _GEN_3276; // @[Sbuffer.scala 160:18]
  wire  _GEN_4925 = wen_12 ? _GEN_4893 : _GEN_3277; // @[Sbuffer.scala 160:18]
  wire  _GEN_4926 = wen_12 ? _GEN_4894 : _GEN_3278; // @[Sbuffer.scala 160:18]
  wire  _GEN_4927 = wen_12 ? _GEN_4895 : _GEN_3279; // @[Sbuffer.scala 160:18]
  wire  _wen_T_55 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_13 = w_valid_s1_0 & _wen_T_55; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4928 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4929 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4930 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4931 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4932 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4933 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4934 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4935 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4936 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4937 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4938 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4939 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4940 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4941 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4942 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4943 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_1_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_4944 = 4'h0 == w_addr_s1_0 | _GEN_3280; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4945 = 4'h1 == w_addr_s1_0 | _GEN_3281; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4946 = 4'h2 == w_addr_s1_0 | _GEN_3282; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4947 = 4'h3 == w_addr_s1_0 | _GEN_3283; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4948 = 4'h4 == w_addr_s1_0 | _GEN_3284; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4949 = 4'h5 == w_addr_s1_0 | _GEN_3285; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4950 = 4'h6 == w_addr_s1_0 | _GEN_3286; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4951 = 4'h7 == w_addr_s1_0 | _GEN_3287; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4952 = 4'h8 == w_addr_s1_0 | _GEN_3288; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4953 = 4'h9 == w_addr_s1_0 | _GEN_3289; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4954 = 4'ha == w_addr_s1_0 | _GEN_3290; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4955 = 4'hb == w_addr_s1_0 | _GEN_3291; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4956 = 4'hc == w_addr_s1_0 | _GEN_3292; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4957 = 4'hd == w_addr_s1_0 | _GEN_3293; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4958 = 4'he == w_addr_s1_0 | _GEN_3294; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_4959 = 4'hf == w_addr_s1_0 | _GEN_3295; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_4960 = wen_13 ? _GEN_4928 : data_0_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4961 = wen_13 ? _GEN_4929 : data_1_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4962 = wen_13 ? _GEN_4930 : data_2_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4963 = wen_13 ? _GEN_4931 : data_3_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4964 = wen_13 ? _GEN_4932 : data_4_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4965 = wen_13 ? _GEN_4933 : data_5_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4966 = wen_13 ? _GEN_4934 : data_6_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4967 = wen_13 ? _GEN_4935 : data_7_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4968 = wen_13 ? _GEN_4936 : data_8_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4969 = wen_13 ? _GEN_4937 : data_9_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4970 = wen_13 ? _GEN_4938 : data_10_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4971 = wen_13 ? _GEN_4939 : data_11_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4972 = wen_13 ? _GEN_4940 : data_12_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4973 = wen_13 ? _GEN_4941 : data_13_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4974 = wen_13 ? _GEN_4942 : data_14_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_4975 = wen_13 ? _GEN_4943 : data_15_1_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_4976 = wen_13 ? _GEN_4944 : _GEN_3280; // @[Sbuffer.scala 160:18]
  wire  _GEN_4977 = wen_13 ? _GEN_4945 : _GEN_3281; // @[Sbuffer.scala 160:18]
  wire  _GEN_4978 = wen_13 ? _GEN_4946 : _GEN_3282; // @[Sbuffer.scala 160:18]
  wire  _GEN_4979 = wen_13 ? _GEN_4947 : _GEN_3283; // @[Sbuffer.scala 160:18]
  wire  _GEN_4980 = wen_13 ? _GEN_4948 : _GEN_3284; // @[Sbuffer.scala 160:18]
  wire  _GEN_4981 = wen_13 ? _GEN_4949 : _GEN_3285; // @[Sbuffer.scala 160:18]
  wire  _GEN_4982 = wen_13 ? _GEN_4950 : _GEN_3286; // @[Sbuffer.scala 160:18]
  wire  _GEN_4983 = wen_13 ? _GEN_4951 : _GEN_3287; // @[Sbuffer.scala 160:18]
  wire  _GEN_4984 = wen_13 ? _GEN_4952 : _GEN_3288; // @[Sbuffer.scala 160:18]
  wire  _GEN_4985 = wen_13 ? _GEN_4953 : _GEN_3289; // @[Sbuffer.scala 160:18]
  wire  _GEN_4986 = wen_13 ? _GEN_4954 : _GEN_3290; // @[Sbuffer.scala 160:18]
  wire  _GEN_4987 = wen_13 ? _GEN_4955 : _GEN_3291; // @[Sbuffer.scala 160:18]
  wire  _GEN_4988 = wen_13 ? _GEN_4956 : _GEN_3292; // @[Sbuffer.scala 160:18]
  wire  _GEN_4989 = wen_13 ? _GEN_4957 : _GEN_3293; // @[Sbuffer.scala 160:18]
  wire  _GEN_4990 = wen_13 ? _GEN_4958 : _GEN_3294; // @[Sbuffer.scala 160:18]
  wire  _GEN_4991 = wen_13 ? _GEN_4959 : _GEN_3295; // @[Sbuffer.scala 160:18]
  wire  _wen_T_59 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_14 = w_valid_s1_0 & _wen_T_59; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_4992 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4993 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4994 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4995 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4996 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4997 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4998 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_4999 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5000 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5001 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5002 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5003 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5004 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5005 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5006 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5007 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_1_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5008 = 4'h0 == w_addr_s1_0 | _GEN_3296; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5009 = 4'h1 == w_addr_s1_0 | _GEN_3297; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5010 = 4'h2 == w_addr_s1_0 | _GEN_3298; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5011 = 4'h3 == w_addr_s1_0 | _GEN_3299; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5012 = 4'h4 == w_addr_s1_0 | _GEN_3300; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5013 = 4'h5 == w_addr_s1_0 | _GEN_3301; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5014 = 4'h6 == w_addr_s1_0 | _GEN_3302; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5015 = 4'h7 == w_addr_s1_0 | _GEN_3303; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5016 = 4'h8 == w_addr_s1_0 | _GEN_3304; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5017 = 4'h9 == w_addr_s1_0 | _GEN_3305; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5018 = 4'ha == w_addr_s1_0 | _GEN_3306; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5019 = 4'hb == w_addr_s1_0 | _GEN_3307; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5020 = 4'hc == w_addr_s1_0 | _GEN_3308; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5021 = 4'hd == w_addr_s1_0 | _GEN_3309; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5022 = 4'he == w_addr_s1_0 | _GEN_3310; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5023 = 4'hf == w_addr_s1_0 | _GEN_3311; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5024 = wen_14 ? _GEN_4992 : data_0_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5025 = wen_14 ? _GEN_4993 : data_1_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5026 = wen_14 ? _GEN_4994 : data_2_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5027 = wen_14 ? _GEN_4995 : data_3_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5028 = wen_14 ? _GEN_4996 : data_4_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5029 = wen_14 ? _GEN_4997 : data_5_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5030 = wen_14 ? _GEN_4998 : data_6_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5031 = wen_14 ? _GEN_4999 : data_7_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5032 = wen_14 ? _GEN_5000 : data_8_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5033 = wen_14 ? _GEN_5001 : data_9_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5034 = wen_14 ? _GEN_5002 : data_10_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5035 = wen_14 ? _GEN_5003 : data_11_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5036 = wen_14 ? _GEN_5004 : data_12_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5037 = wen_14 ? _GEN_5005 : data_13_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5038 = wen_14 ? _GEN_5006 : data_14_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5039 = wen_14 ? _GEN_5007 : data_15_1_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5040 = wen_14 ? _GEN_5008 : _GEN_3296; // @[Sbuffer.scala 160:18]
  wire  _GEN_5041 = wen_14 ? _GEN_5009 : _GEN_3297; // @[Sbuffer.scala 160:18]
  wire  _GEN_5042 = wen_14 ? _GEN_5010 : _GEN_3298; // @[Sbuffer.scala 160:18]
  wire  _GEN_5043 = wen_14 ? _GEN_5011 : _GEN_3299; // @[Sbuffer.scala 160:18]
  wire  _GEN_5044 = wen_14 ? _GEN_5012 : _GEN_3300; // @[Sbuffer.scala 160:18]
  wire  _GEN_5045 = wen_14 ? _GEN_5013 : _GEN_3301; // @[Sbuffer.scala 160:18]
  wire  _GEN_5046 = wen_14 ? _GEN_5014 : _GEN_3302; // @[Sbuffer.scala 160:18]
  wire  _GEN_5047 = wen_14 ? _GEN_5015 : _GEN_3303; // @[Sbuffer.scala 160:18]
  wire  _GEN_5048 = wen_14 ? _GEN_5016 : _GEN_3304; // @[Sbuffer.scala 160:18]
  wire  _GEN_5049 = wen_14 ? _GEN_5017 : _GEN_3305; // @[Sbuffer.scala 160:18]
  wire  _GEN_5050 = wen_14 ? _GEN_5018 : _GEN_3306; // @[Sbuffer.scala 160:18]
  wire  _GEN_5051 = wen_14 ? _GEN_5019 : _GEN_3307; // @[Sbuffer.scala 160:18]
  wire  _GEN_5052 = wen_14 ? _GEN_5020 : _GEN_3308; // @[Sbuffer.scala 160:18]
  wire  _GEN_5053 = wen_14 ? _GEN_5021 : _GEN_3309; // @[Sbuffer.scala 160:18]
  wire  _GEN_5054 = wen_14 ? _GEN_5022 : _GEN_3310; // @[Sbuffer.scala 160:18]
  wire  _GEN_5055 = wen_14 ? _GEN_5023 : _GEN_3311; // @[Sbuffer.scala 160:18]
  wire  _wen_T_63 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h1 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_15 = w_valid_s1_0 & _wen_T_63; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5056 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5057 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5058 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5059 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5060 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5061 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5062 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5063 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5064 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5065 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5066 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5067 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5068 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5069 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5070 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5071 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_1_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5072 = 4'h0 == w_addr_s1_0 | _GEN_3312; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5073 = 4'h1 == w_addr_s1_0 | _GEN_3313; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5074 = 4'h2 == w_addr_s1_0 | _GEN_3314; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5075 = 4'h3 == w_addr_s1_0 | _GEN_3315; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5076 = 4'h4 == w_addr_s1_0 | _GEN_3316; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5077 = 4'h5 == w_addr_s1_0 | _GEN_3317; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5078 = 4'h6 == w_addr_s1_0 | _GEN_3318; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5079 = 4'h7 == w_addr_s1_0 | _GEN_3319; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5080 = 4'h8 == w_addr_s1_0 | _GEN_3320; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5081 = 4'h9 == w_addr_s1_0 | _GEN_3321; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5082 = 4'ha == w_addr_s1_0 | _GEN_3322; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5083 = 4'hb == w_addr_s1_0 | _GEN_3323; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5084 = 4'hc == w_addr_s1_0 | _GEN_3324; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5085 = 4'hd == w_addr_s1_0 | _GEN_3325; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5086 = 4'he == w_addr_s1_0 | _GEN_3326; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5087 = 4'hf == w_addr_s1_0 | _GEN_3327; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5088 = wen_15 ? _GEN_5056 : data_0_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5089 = wen_15 ? _GEN_5057 : data_1_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5090 = wen_15 ? _GEN_5058 : data_2_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5091 = wen_15 ? _GEN_5059 : data_3_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5092 = wen_15 ? _GEN_5060 : data_4_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5093 = wen_15 ? _GEN_5061 : data_5_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5094 = wen_15 ? _GEN_5062 : data_6_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5095 = wen_15 ? _GEN_5063 : data_7_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5096 = wen_15 ? _GEN_5064 : data_8_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5097 = wen_15 ? _GEN_5065 : data_9_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5098 = wen_15 ? _GEN_5066 : data_10_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5099 = wen_15 ? _GEN_5067 : data_11_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5100 = wen_15 ? _GEN_5068 : data_12_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5101 = wen_15 ? _GEN_5069 : data_13_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5102 = wen_15 ? _GEN_5070 : data_14_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5103 = wen_15 ? _GEN_5071 : data_15_1_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5104 = wen_15 ? _GEN_5072 : _GEN_3312; // @[Sbuffer.scala 160:18]
  wire  _GEN_5105 = wen_15 ? _GEN_5073 : _GEN_3313; // @[Sbuffer.scala 160:18]
  wire  _GEN_5106 = wen_15 ? _GEN_5074 : _GEN_3314; // @[Sbuffer.scala 160:18]
  wire  _GEN_5107 = wen_15 ? _GEN_5075 : _GEN_3315; // @[Sbuffer.scala 160:18]
  wire  _GEN_5108 = wen_15 ? _GEN_5076 : _GEN_3316; // @[Sbuffer.scala 160:18]
  wire  _GEN_5109 = wen_15 ? _GEN_5077 : _GEN_3317; // @[Sbuffer.scala 160:18]
  wire  _GEN_5110 = wen_15 ? _GEN_5078 : _GEN_3318; // @[Sbuffer.scala 160:18]
  wire  _GEN_5111 = wen_15 ? _GEN_5079 : _GEN_3319; // @[Sbuffer.scala 160:18]
  wire  _GEN_5112 = wen_15 ? _GEN_5080 : _GEN_3320; // @[Sbuffer.scala 160:18]
  wire  _GEN_5113 = wen_15 ? _GEN_5081 : _GEN_3321; // @[Sbuffer.scala 160:18]
  wire  _GEN_5114 = wen_15 ? _GEN_5082 : _GEN_3322; // @[Sbuffer.scala 160:18]
  wire  _GEN_5115 = wen_15 ? _GEN_5083 : _GEN_3323; // @[Sbuffer.scala 160:18]
  wire  _GEN_5116 = wen_15 ? _GEN_5084 : _GEN_3324; // @[Sbuffer.scala 160:18]
  wire  _GEN_5117 = wen_15 ? _GEN_5085 : _GEN_3325; // @[Sbuffer.scala 160:18]
  wire  _GEN_5118 = wen_15 ? _GEN_5086 : _GEN_3326; // @[Sbuffer.scala 160:18]
  wire  _GEN_5119 = wen_15 ? _GEN_5087 : _GEN_3327; // @[Sbuffer.scala 160:18]
  wire  _wen_T_67 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_16 = w_valid_s1_0 & _wen_T_67; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5120 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5121 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5122 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5123 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5124 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5125 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5126 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5127 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5128 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5129 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5130 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5131 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5132 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5133 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5134 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5135 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_2_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5136 = 4'h0 == w_addr_s1_0 | _GEN_3328; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5137 = 4'h1 == w_addr_s1_0 | _GEN_3329; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5138 = 4'h2 == w_addr_s1_0 | _GEN_3330; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5139 = 4'h3 == w_addr_s1_0 | _GEN_3331; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5140 = 4'h4 == w_addr_s1_0 | _GEN_3332; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5141 = 4'h5 == w_addr_s1_0 | _GEN_3333; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5142 = 4'h6 == w_addr_s1_0 | _GEN_3334; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5143 = 4'h7 == w_addr_s1_0 | _GEN_3335; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5144 = 4'h8 == w_addr_s1_0 | _GEN_3336; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5145 = 4'h9 == w_addr_s1_0 | _GEN_3337; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5146 = 4'ha == w_addr_s1_0 | _GEN_3338; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5147 = 4'hb == w_addr_s1_0 | _GEN_3339; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5148 = 4'hc == w_addr_s1_0 | _GEN_3340; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5149 = 4'hd == w_addr_s1_0 | _GEN_3341; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5150 = 4'he == w_addr_s1_0 | _GEN_3342; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5151 = 4'hf == w_addr_s1_0 | _GEN_3343; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5152 = wen_16 ? _GEN_5120 : data_0_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5153 = wen_16 ? _GEN_5121 : data_1_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5154 = wen_16 ? _GEN_5122 : data_2_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5155 = wen_16 ? _GEN_5123 : data_3_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5156 = wen_16 ? _GEN_5124 : data_4_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5157 = wen_16 ? _GEN_5125 : data_5_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5158 = wen_16 ? _GEN_5126 : data_6_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5159 = wen_16 ? _GEN_5127 : data_7_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5160 = wen_16 ? _GEN_5128 : data_8_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5161 = wen_16 ? _GEN_5129 : data_9_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5162 = wen_16 ? _GEN_5130 : data_10_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5163 = wen_16 ? _GEN_5131 : data_11_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5164 = wen_16 ? _GEN_5132 : data_12_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5165 = wen_16 ? _GEN_5133 : data_13_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5166 = wen_16 ? _GEN_5134 : data_14_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5167 = wen_16 ? _GEN_5135 : data_15_2_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5168 = wen_16 ? _GEN_5136 : _GEN_3328; // @[Sbuffer.scala 160:18]
  wire  _GEN_5169 = wen_16 ? _GEN_5137 : _GEN_3329; // @[Sbuffer.scala 160:18]
  wire  _GEN_5170 = wen_16 ? _GEN_5138 : _GEN_3330; // @[Sbuffer.scala 160:18]
  wire  _GEN_5171 = wen_16 ? _GEN_5139 : _GEN_3331; // @[Sbuffer.scala 160:18]
  wire  _GEN_5172 = wen_16 ? _GEN_5140 : _GEN_3332; // @[Sbuffer.scala 160:18]
  wire  _GEN_5173 = wen_16 ? _GEN_5141 : _GEN_3333; // @[Sbuffer.scala 160:18]
  wire  _GEN_5174 = wen_16 ? _GEN_5142 : _GEN_3334; // @[Sbuffer.scala 160:18]
  wire  _GEN_5175 = wen_16 ? _GEN_5143 : _GEN_3335; // @[Sbuffer.scala 160:18]
  wire  _GEN_5176 = wen_16 ? _GEN_5144 : _GEN_3336; // @[Sbuffer.scala 160:18]
  wire  _GEN_5177 = wen_16 ? _GEN_5145 : _GEN_3337; // @[Sbuffer.scala 160:18]
  wire  _GEN_5178 = wen_16 ? _GEN_5146 : _GEN_3338; // @[Sbuffer.scala 160:18]
  wire  _GEN_5179 = wen_16 ? _GEN_5147 : _GEN_3339; // @[Sbuffer.scala 160:18]
  wire  _GEN_5180 = wen_16 ? _GEN_5148 : _GEN_3340; // @[Sbuffer.scala 160:18]
  wire  _GEN_5181 = wen_16 ? _GEN_5149 : _GEN_3341; // @[Sbuffer.scala 160:18]
  wire  _GEN_5182 = wen_16 ? _GEN_5150 : _GEN_3342; // @[Sbuffer.scala 160:18]
  wire  _GEN_5183 = wen_16 ? _GEN_5151 : _GEN_3343; // @[Sbuffer.scala 160:18]
  wire  _wen_T_71 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_17 = w_valid_s1_0 & _wen_T_71; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5184 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5185 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5186 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5187 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5188 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5189 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5190 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5191 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5192 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5193 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5194 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5195 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5196 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5197 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5198 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5199 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_2_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5200 = 4'h0 == w_addr_s1_0 | _GEN_3344; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5201 = 4'h1 == w_addr_s1_0 | _GEN_3345; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5202 = 4'h2 == w_addr_s1_0 | _GEN_3346; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5203 = 4'h3 == w_addr_s1_0 | _GEN_3347; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5204 = 4'h4 == w_addr_s1_0 | _GEN_3348; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5205 = 4'h5 == w_addr_s1_0 | _GEN_3349; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5206 = 4'h6 == w_addr_s1_0 | _GEN_3350; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5207 = 4'h7 == w_addr_s1_0 | _GEN_3351; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5208 = 4'h8 == w_addr_s1_0 | _GEN_3352; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5209 = 4'h9 == w_addr_s1_0 | _GEN_3353; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5210 = 4'ha == w_addr_s1_0 | _GEN_3354; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5211 = 4'hb == w_addr_s1_0 | _GEN_3355; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5212 = 4'hc == w_addr_s1_0 | _GEN_3356; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5213 = 4'hd == w_addr_s1_0 | _GEN_3357; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5214 = 4'he == w_addr_s1_0 | _GEN_3358; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5215 = 4'hf == w_addr_s1_0 | _GEN_3359; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5216 = wen_17 ? _GEN_5184 : data_0_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5217 = wen_17 ? _GEN_5185 : data_1_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5218 = wen_17 ? _GEN_5186 : data_2_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5219 = wen_17 ? _GEN_5187 : data_3_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5220 = wen_17 ? _GEN_5188 : data_4_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5221 = wen_17 ? _GEN_5189 : data_5_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5222 = wen_17 ? _GEN_5190 : data_6_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5223 = wen_17 ? _GEN_5191 : data_7_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5224 = wen_17 ? _GEN_5192 : data_8_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5225 = wen_17 ? _GEN_5193 : data_9_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5226 = wen_17 ? _GEN_5194 : data_10_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5227 = wen_17 ? _GEN_5195 : data_11_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5228 = wen_17 ? _GEN_5196 : data_12_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5229 = wen_17 ? _GEN_5197 : data_13_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5230 = wen_17 ? _GEN_5198 : data_14_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5231 = wen_17 ? _GEN_5199 : data_15_2_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5232 = wen_17 ? _GEN_5200 : _GEN_3344; // @[Sbuffer.scala 160:18]
  wire  _GEN_5233 = wen_17 ? _GEN_5201 : _GEN_3345; // @[Sbuffer.scala 160:18]
  wire  _GEN_5234 = wen_17 ? _GEN_5202 : _GEN_3346; // @[Sbuffer.scala 160:18]
  wire  _GEN_5235 = wen_17 ? _GEN_5203 : _GEN_3347; // @[Sbuffer.scala 160:18]
  wire  _GEN_5236 = wen_17 ? _GEN_5204 : _GEN_3348; // @[Sbuffer.scala 160:18]
  wire  _GEN_5237 = wen_17 ? _GEN_5205 : _GEN_3349; // @[Sbuffer.scala 160:18]
  wire  _GEN_5238 = wen_17 ? _GEN_5206 : _GEN_3350; // @[Sbuffer.scala 160:18]
  wire  _GEN_5239 = wen_17 ? _GEN_5207 : _GEN_3351; // @[Sbuffer.scala 160:18]
  wire  _GEN_5240 = wen_17 ? _GEN_5208 : _GEN_3352; // @[Sbuffer.scala 160:18]
  wire  _GEN_5241 = wen_17 ? _GEN_5209 : _GEN_3353; // @[Sbuffer.scala 160:18]
  wire  _GEN_5242 = wen_17 ? _GEN_5210 : _GEN_3354; // @[Sbuffer.scala 160:18]
  wire  _GEN_5243 = wen_17 ? _GEN_5211 : _GEN_3355; // @[Sbuffer.scala 160:18]
  wire  _GEN_5244 = wen_17 ? _GEN_5212 : _GEN_3356; // @[Sbuffer.scala 160:18]
  wire  _GEN_5245 = wen_17 ? _GEN_5213 : _GEN_3357; // @[Sbuffer.scala 160:18]
  wire  _GEN_5246 = wen_17 ? _GEN_5214 : _GEN_3358; // @[Sbuffer.scala 160:18]
  wire  _GEN_5247 = wen_17 ? _GEN_5215 : _GEN_3359; // @[Sbuffer.scala 160:18]
  wire  _wen_T_75 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_18 = w_valid_s1_0 & _wen_T_75; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5248 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5249 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5250 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5251 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5252 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5253 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5254 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5255 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5256 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5257 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5258 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5259 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5260 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5261 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5262 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5263 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_2_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5264 = 4'h0 == w_addr_s1_0 | _GEN_3360; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5265 = 4'h1 == w_addr_s1_0 | _GEN_3361; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5266 = 4'h2 == w_addr_s1_0 | _GEN_3362; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5267 = 4'h3 == w_addr_s1_0 | _GEN_3363; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5268 = 4'h4 == w_addr_s1_0 | _GEN_3364; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5269 = 4'h5 == w_addr_s1_0 | _GEN_3365; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5270 = 4'h6 == w_addr_s1_0 | _GEN_3366; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5271 = 4'h7 == w_addr_s1_0 | _GEN_3367; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5272 = 4'h8 == w_addr_s1_0 | _GEN_3368; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5273 = 4'h9 == w_addr_s1_0 | _GEN_3369; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5274 = 4'ha == w_addr_s1_0 | _GEN_3370; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5275 = 4'hb == w_addr_s1_0 | _GEN_3371; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5276 = 4'hc == w_addr_s1_0 | _GEN_3372; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5277 = 4'hd == w_addr_s1_0 | _GEN_3373; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5278 = 4'he == w_addr_s1_0 | _GEN_3374; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5279 = 4'hf == w_addr_s1_0 | _GEN_3375; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5280 = wen_18 ? _GEN_5248 : data_0_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5281 = wen_18 ? _GEN_5249 : data_1_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5282 = wen_18 ? _GEN_5250 : data_2_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5283 = wen_18 ? _GEN_5251 : data_3_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5284 = wen_18 ? _GEN_5252 : data_4_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5285 = wen_18 ? _GEN_5253 : data_5_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5286 = wen_18 ? _GEN_5254 : data_6_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5287 = wen_18 ? _GEN_5255 : data_7_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5288 = wen_18 ? _GEN_5256 : data_8_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5289 = wen_18 ? _GEN_5257 : data_9_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5290 = wen_18 ? _GEN_5258 : data_10_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5291 = wen_18 ? _GEN_5259 : data_11_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5292 = wen_18 ? _GEN_5260 : data_12_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5293 = wen_18 ? _GEN_5261 : data_13_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5294 = wen_18 ? _GEN_5262 : data_14_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5295 = wen_18 ? _GEN_5263 : data_15_2_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5296 = wen_18 ? _GEN_5264 : _GEN_3360; // @[Sbuffer.scala 160:18]
  wire  _GEN_5297 = wen_18 ? _GEN_5265 : _GEN_3361; // @[Sbuffer.scala 160:18]
  wire  _GEN_5298 = wen_18 ? _GEN_5266 : _GEN_3362; // @[Sbuffer.scala 160:18]
  wire  _GEN_5299 = wen_18 ? _GEN_5267 : _GEN_3363; // @[Sbuffer.scala 160:18]
  wire  _GEN_5300 = wen_18 ? _GEN_5268 : _GEN_3364; // @[Sbuffer.scala 160:18]
  wire  _GEN_5301 = wen_18 ? _GEN_5269 : _GEN_3365; // @[Sbuffer.scala 160:18]
  wire  _GEN_5302 = wen_18 ? _GEN_5270 : _GEN_3366; // @[Sbuffer.scala 160:18]
  wire  _GEN_5303 = wen_18 ? _GEN_5271 : _GEN_3367; // @[Sbuffer.scala 160:18]
  wire  _GEN_5304 = wen_18 ? _GEN_5272 : _GEN_3368; // @[Sbuffer.scala 160:18]
  wire  _GEN_5305 = wen_18 ? _GEN_5273 : _GEN_3369; // @[Sbuffer.scala 160:18]
  wire  _GEN_5306 = wen_18 ? _GEN_5274 : _GEN_3370; // @[Sbuffer.scala 160:18]
  wire  _GEN_5307 = wen_18 ? _GEN_5275 : _GEN_3371; // @[Sbuffer.scala 160:18]
  wire  _GEN_5308 = wen_18 ? _GEN_5276 : _GEN_3372; // @[Sbuffer.scala 160:18]
  wire  _GEN_5309 = wen_18 ? _GEN_5277 : _GEN_3373; // @[Sbuffer.scala 160:18]
  wire  _GEN_5310 = wen_18 ? _GEN_5278 : _GEN_3374; // @[Sbuffer.scala 160:18]
  wire  _GEN_5311 = wen_18 ? _GEN_5279 : _GEN_3375; // @[Sbuffer.scala 160:18]
  wire  _wen_T_79 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_19 = w_valid_s1_0 & _wen_T_79; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5312 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5313 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5314 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5315 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5316 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5317 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5318 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5319 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5320 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5321 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5322 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5323 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5324 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5325 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5326 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5327 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_2_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5328 = 4'h0 == w_addr_s1_0 | _GEN_3376; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5329 = 4'h1 == w_addr_s1_0 | _GEN_3377; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5330 = 4'h2 == w_addr_s1_0 | _GEN_3378; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5331 = 4'h3 == w_addr_s1_0 | _GEN_3379; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5332 = 4'h4 == w_addr_s1_0 | _GEN_3380; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5333 = 4'h5 == w_addr_s1_0 | _GEN_3381; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5334 = 4'h6 == w_addr_s1_0 | _GEN_3382; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5335 = 4'h7 == w_addr_s1_0 | _GEN_3383; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5336 = 4'h8 == w_addr_s1_0 | _GEN_3384; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5337 = 4'h9 == w_addr_s1_0 | _GEN_3385; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5338 = 4'ha == w_addr_s1_0 | _GEN_3386; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5339 = 4'hb == w_addr_s1_0 | _GEN_3387; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5340 = 4'hc == w_addr_s1_0 | _GEN_3388; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5341 = 4'hd == w_addr_s1_0 | _GEN_3389; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5342 = 4'he == w_addr_s1_0 | _GEN_3390; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5343 = 4'hf == w_addr_s1_0 | _GEN_3391; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5344 = wen_19 ? _GEN_5312 : data_0_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5345 = wen_19 ? _GEN_5313 : data_1_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5346 = wen_19 ? _GEN_5314 : data_2_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5347 = wen_19 ? _GEN_5315 : data_3_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5348 = wen_19 ? _GEN_5316 : data_4_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5349 = wen_19 ? _GEN_5317 : data_5_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5350 = wen_19 ? _GEN_5318 : data_6_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5351 = wen_19 ? _GEN_5319 : data_7_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5352 = wen_19 ? _GEN_5320 : data_8_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5353 = wen_19 ? _GEN_5321 : data_9_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5354 = wen_19 ? _GEN_5322 : data_10_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5355 = wen_19 ? _GEN_5323 : data_11_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5356 = wen_19 ? _GEN_5324 : data_12_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5357 = wen_19 ? _GEN_5325 : data_13_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5358 = wen_19 ? _GEN_5326 : data_14_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5359 = wen_19 ? _GEN_5327 : data_15_2_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5360 = wen_19 ? _GEN_5328 : _GEN_3376; // @[Sbuffer.scala 160:18]
  wire  _GEN_5361 = wen_19 ? _GEN_5329 : _GEN_3377; // @[Sbuffer.scala 160:18]
  wire  _GEN_5362 = wen_19 ? _GEN_5330 : _GEN_3378; // @[Sbuffer.scala 160:18]
  wire  _GEN_5363 = wen_19 ? _GEN_5331 : _GEN_3379; // @[Sbuffer.scala 160:18]
  wire  _GEN_5364 = wen_19 ? _GEN_5332 : _GEN_3380; // @[Sbuffer.scala 160:18]
  wire  _GEN_5365 = wen_19 ? _GEN_5333 : _GEN_3381; // @[Sbuffer.scala 160:18]
  wire  _GEN_5366 = wen_19 ? _GEN_5334 : _GEN_3382; // @[Sbuffer.scala 160:18]
  wire  _GEN_5367 = wen_19 ? _GEN_5335 : _GEN_3383; // @[Sbuffer.scala 160:18]
  wire  _GEN_5368 = wen_19 ? _GEN_5336 : _GEN_3384; // @[Sbuffer.scala 160:18]
  wire  _GEN_5369 = wen_19 ? _GEN_5337 : _GEN_3385; // @[Sbuffer.scala 160:18]
  wire  _GEN_5370 = wen_19 ? _GEN_5338 : _GEN_3386; // @[Sbuffer.scala 160:18]
  wire  _GEN_5371 = wen_19 ? _GEN_5339 : _GEN_3387; // @[Sbuffer.scala 160:18]
  wire  _GEN_5372 = wen_19 ? _GEN_5340 : _GEN_3388; // @[Sbuffer.scala 160:18]
  wire  _GEN_5373 = wen_19 ? _GEN_5341 : _GEN_3389; // @[Sbuffer.scala 160:18]
  wire  _GEN_5374 = wen_19 ? _GEN_5342 : _GEN_3390; // @[Sbuffer.scala 160:18]
  wire  _GEN_5375 = wen_19 ? _GEN_5343 : _GEN_3391; // @[Sbuffer.scala 160:18]
  wire  _wen_T_83 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_20 = w_valid_s1_0 & _wen_T_83; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5376 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5377 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5378 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5379 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5380 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5381 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5382 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5383 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5384 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5385 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5386 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5387 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5388 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5389 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5390 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5391 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_2_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5392 = 4'h0 == w_addr_s1_0 | _GEN_3392; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5393 = 4'h1 == w_addr_s1_0 | _GEN_3393; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5394 = 4'h2 == w_addr_s1_0 | _GEN_3394; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5395 = 4'h3 == w_addr_s1_0 | _GEN_3395; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5396 = 4'h4 == w_addr_s1_0 | _GEN_3396; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5397 = 4'h5 == w_addr_s1_0 | _GEN_3397; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5398 = 4'h6 == w_addr_s1_0 | _GEN_3398; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5399 = 4'h7 == w_addr_s1_0 | _GEN_3399; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5400 = 4'h8 == w_addr_s1_0 | _GEN_3400; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5401 = 4'h9 == w_addr_s1_0 | _GEN_3401; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5402 = 4'ha == w_addr_s1_0 | _GEN_3402; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5403 = 4'hb == w_addr_s1_0 | _GEN_3403; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5404 = 4'hc == w_addr_s1_0 | _GEN_3404; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5405 = 4'hd == w_addr_s1_0 | _GEN_3405; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5406 = 4'he == w_addr_s1_0 | _GEN_3406; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5407 = 4'hf == w_addr_s1_0 | _GEN_3407; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5408 = wen_20 ? _GEN_5376 : data_0_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5409 = wen_20 ? _GEN_5377 : data_1_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5410 = wen_20 ? _GEN_5378 : data_2_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5411 = wen_20 ? _GEN_5379 : data_3_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5412 = wen_20 ? _GEN_5380 : data_4_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5413 = wen_20 ? _GEN_5381 : data_5_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5414 = wen_20 ? _GEN_5382 : data_6_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5415 = wen_20 ? _GEN_5383 : data_7_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5416 = wen_20 ? _GEN_5384 : data_8_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5417 = wen_20 ? _GEN_5385 : data_9_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5418 = wen_20 ? _GEN_5386 : data_10_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5419 = wen_20 ? _GEN_5387 : data_11_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5420 = wen_20 ? _GEN_5388 : data_12_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5421 = wen_20 ? _GEN_5389 : data_13_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5422 = wen_20 ? _GEN_5390 : data_14_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5423 = wen_20 ? _GEN_5391 : data_15_2_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5424 = wen_20 ? _GEN_5392 : _GEN_3392; // @[Sbuffer.scala 160:18]
  wire  _GEN_5425 = wen_20 ? _GEN_5393 : _GEN_3393; // @[Sbuffer.scala 160:18]
  wire  _GEN_5426 = wen_20 ? _GEN_5394 : _GEN_3394; // @[Sbuffer.scala 160:18]
  wire  _GEN_5427 = wen_20 ? _GEN_5395 : _GEN_3395; // @[Sbuffer.scala 160:18]
  wire  _GEN_5428 = wen_20 ? _GEN_5396 : _GEN_3396; // @[Sbuffer.scala 160:18]
  wire  _GEN_5429 = wen_20 ? _GEN_5397 : _GEN_3397; // @[Sbuffer.scala 160:18]
  wire  _GEN_5430 = wen_20 ? _GEN_5398 : _GEN_3398; // @[Sbuffer.scala 160:18]
  wire  _GEN_5431 = wen_20 ? _GEN_5399 : _GEN_3399; // @[Sbuffer.scala 160:18]
  wire  _GEN_5432 = wen_20 ? _GEN_5400 : _GEN_3400; // @[Sbuffer.scala 160:18]
  wire  _GEN_5433 = wen_20 ? _GEN_5401 : _GEN_3401; // @[Sbuffer.scala 160:18]
  wire  _GEN_5434 = wen_20 ? _GEN_5402 : _GEN_3402; // @[Sbuffer.scala 160:18]
  wire  _GEN_5435 = wen_20 ? _GEN_5403 : _GEN_3403; // @[Sbuffer.scala 160:18]
  wire  _GEN_5436 = wen_20 ? _GEN_5404 : _GEN_3404; // @[Sbuffer.scala 160:18]
  wire  _GEN_5437 = wen_20 ? _GEN_5405 : _GEN_3405; // @[Sbuffer.scala 160:18]
  wire  _GEN_5438 = wen_20 ? _GEN_5406 : _GEN_3406; // @[Sbuffer.scala 160:18]
  wire  _GEN_5439 = wen_20 ? _GEN_5407 : _GEN_3407; // @[Sbuffer.scala 160:18]
  wire  _wen_T_87 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_21 = w_valid_s1_0 & _wen_T_87; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5440 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5441 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5442 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5443 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5444 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5445 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5446 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5447 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5448 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5449 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5450 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5451 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5452 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5453 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5454 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5455 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_2_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5456 = 4'h0 == w_addr_s1_0 | _GEN_3408; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5457 = 4'h1 == w_addr_s1_0 | _GEN_3409; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5458 = 4'h2 == w_addr_s1_0 | _GEN_3410; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5459 = 4'h3 == w_addr_s1_0 | _GEN_3411; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5460 = 4'h4 == w_addr_s1_0 | _GEN_3412; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5461 = 4'h5 == w_addr_s1_0 | _GEN_3413; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5462 = 4'h6 == w_addr_s1_0 | _GEN_3414; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5463 = 4'h7 == w_addr_s1_0 | _GEN_3415; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5464 = 4'h8 == w_addr_s1_0 | _GEN_3416; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5465 = 4'h9 == w_addr_s1_0 | _GEN_3417; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5466 = 4'ha == w_addr_s1_0 | _GEN_3418; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5467 = 4'hb == w_addr_s1_0 | _GEN_3419; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5468 = 4'hc == w_addr_s1_0 | _GEN_3420; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5469 = 4'hd == w_addr_s1_0 | _GEN_3421; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5470 = 4'he == w_addr_s1_0 | _GEN_3422; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5471 = 4'hf == w_addr_s1_0 | _GEN_3423; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5472 = wen_21 ? _GEN_5440 : data_0_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5473 = wen_21 ? _GEN_5441 : data_1_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5474 = wen_21 ? _GEN_5442 : data_2_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5475 = wen_21 ? _GEN_5443 : data_3_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5476 = wen_21 ? _GEN_5444 : data_4_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5477 = wen_21 ? _GEN_5445 : data_5_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5478 = wen_21 ? _GEN_5446 : data_6_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5479 = wen_21 ? _GEN_5447 : data_7_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5480 = wen_21 ? _GEN_5448 : data_8_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5481 = wen_21 ? _GEN_5449 : data_9_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5482 = wen_21 ? _GEN_5450 : data_10_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5483 = wen_21 ? _GEN_5451 : data_11_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5484 = wen_21 ? _GEN_5452 : data_12_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5485 = wen_21 ? _GEN_5453 : data_13_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5486 = wen_21 ? _GEN_5454 : data_14_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5487 = wen_21 ? _GEN_5455 : data_15_2_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5488 = wen_21 ? _GEN_5456 : _GEN_3408; // @[Sbuffer.scala 160:18]
  wire  _GEN_5489 = wen_21 ? _GEN_5457 : _GEN_3409; // @[Sbuffer.scala 160:18]
  wire  _GEN_5490 = wen_21 ? _GEN_5458 : _GEN_3410; // @[Sbuffer.scala 160:18]
  wire  _GEN_5491 = wen_21 ? _GEN_5459 : _GEN_3411; // @[Sbuffer.scala 160:18]
  wire  _GEN_5492 = wen_21 ? _GEN_5460 : _GEN_3412; // @[Sbuffer.scala 160:18]
  wire  _GEN_5493 = wen_21 ? _GEN_5461 : _GEN_3413; // @[Sbuffer.scala 160:18]
  wire  _GEN_5494 = wen_21 ? _GEN_5462 : _GEN_3414; // @[Sbuffer.scala 160:18]
  wire  _GEN_5495 = wen_21 ? _GEN_5463 : _GEN_3415; // @[Sbuffer.scala 160:18]
  wire  _GEN_5496 = wen_21 ? _GEN_5464 : _GEN_3416; // @[Sbuffer.scala 160:18]
  wire  _GEN_5497 = wen_21 ? _GEN_5465 : _GEN_3417; // @[Sbuffer.scala 160:18]
  wire  _GEN_5498 = wen_21 ? _GEN_5466 : _GEN_3418; // @[Sbuffer.scala 160:18]
  wire  _GEN_5499 = wen_21 ? _GEN_5467 : _GEN_3419; // @[Sbuffer.scala 160:18]
  wire  _GEN_5500 = wen_21 ? _GEN_5468 : _GEN_3420; // @[Sbuffer.scala 160:18]
  wire  _GEN_5501 = wen_21 ? _GEN_5469 : _GEN_3421; // @[Sbuffer.scala 160:18]
  wire  _GEN_5502 = wen_21 ? _GEN_5470 : _GEN_3422; // @[Sbuffer.scala 160:18]
  wire  _GEN_5503 = wen_21 ? _GEN_5471 : _GEN_3423; // @[Sbuffer.scala 160:18]
  wire  _wen_T_91 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_22 = w_valid_s1_0 & _wen_T_91; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5504 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5505 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5506 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5507 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5508 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5509 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5510 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5511 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5512 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5513 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5514 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5515 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5516 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5517 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5518 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5519 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_2_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5520 = 4'h0 == w_addr_s1_0 | _GEN_3424; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5521 = 4'h1 == w_addr_s1_0 | _GEN_3425; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5522 = 4'h2 == w_addr_s1_0 | _GEN_3426; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5523 = 4'h3 == w_addr_s1_0 | _GEN_3427; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5524 = 4'h4 == w_addr_s1_0 | _GEN_3428; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5525 = 4'h5 == w_addr_s1_0 | _GEN_3429; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5526 = 4'h6 == w_addr_s1_0 | _GEN_3430; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5527 = 4'h7 == w_addr_s1_0 | _GEN_3431; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5528 = 4'h8 == w_addr_s1_0 | _GEN_3432; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5529 = 4'h9 == w_addr_s1_0 | _GEN_3433; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5530 = 4'ha == w_addr_s1_0 | _GEN_3434; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5531 = 4'hb == w_addr_s1_0 | _GEN_3435; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5532 = 4'hc == w_addr_s1_0 | _GEN_3436; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5533 = 4'hd == w_addr_s1_0 | _GEN_3437; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5534 = 4'he == w_addr_s1_0 | _GEN_3438; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5535 = 4'hf == w_addr_s1_0 | _GEN_3439; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5536 = wen_22 ? _GEN_5504 : data_0_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5537 = wen_22 ? _GEN_5505 : data_1_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5538 = wen_22 ? _GEN_5506 : data_2_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5539 = wen_22 ? _GEN_5507 : data_3_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5540 = wen_22 ? _GEN_5508 : data_4_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5541 = wen_22 ? _GEN_5509 : data_5_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5542 = wen_22 ? _GEN_5510 : data_6_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5543 = wen_22 ? _GEN_5511 : data_7_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5544 = wen_22 ? _GEN_5512 : data_8_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5545 = wen_22 ? _GEN_5513 : data_9_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5546 = wen_22 ? _GEN_5514 : data_10_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5547 = wen_22 ? _GEN_5515 : data_11_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5548 = wen_22 ? _GEN_5516 : data_12_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5549 = wen_22 ? _GEN_5517 : data_13_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5550 = wen_22 ? _GEN_5518 : data_14_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5551 = wen_22 ? _GEN_5519 : data_15_2_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5552 = wen_22 ? _GEN_5520 : _GEN_3424; // @[Sbuffer.scala 160:18]
  wire  _GEN_5553 = wen_22 ? _GEN_5521 : _GEN_3425; // @[Sbuffer.scala 160:18]
  wire  _GEN_5554 = wen_22 ? _GEN_5522 : _GEN_3426; // @[Sbuffer.scala 160:18]
  wire  _GEN_5555 = wen_22 ? _GEN_5523 : _GEN_3427; // @[Sbuffer.scala 160:18]
  wire  _GEN_5556 = wen_22 ? _GEN_5524 : _GEN_3428; // @[Sbuffer.scala 160:18]
  wire  _GEN_5557 = wen_22 ? _GEN_5525 : _GEN_3429; // @[Sbuffer.scala 160:18]
  wire  _GEN_5558 = wen_22 ? _GEN_5526 : _GEN_3430; // @[Sbuffer.scala 160:18]
  wire  _GEN_5559 = wen_22 ? _GEN_5527 : _GEN_3431; // @[Sbuffer.scala 160:18]
  wire  _GEN_5560 = wen_22 ? _GEN_5528 : _GEN_3432; // @[Sbuffer.scala 160:18]
  wire  _GEN_5561 = wen_22 ? _GEN_5529 : _GEN_3433; // @[Sbuffer.scala 160:18]
  wire  _GEN_5562 = wen_22 ? _GEN_5530 : _GEN_3434; // @[Sbuffer.scala 160:18]
  wire  _GEN_5563 = wen_22 ? _GEN_5531 : _GEN_3435; // @[Sbuffer.scala 160:18]
  wire  _GEN_5564 = wen_22 ? _GEN_5532 : _GEN_3436; // @[Sbuffer.scala 160:18]
  wire  _GEN_5565 = wen_22 ? _GEN_5533 : _GEN_3437; // @[Sbuffer.scala 160:18]
  wire  _GEN_5566 = wen_22 ? _GEN_5534 : _GEN_3438; // @[Sbuffer.scala 160:18]
  wire  _GEN_5567 = wen_22 ? _GEN_5535 : _GEN_3439; // @[Sbuffer.scala 160:18]
  wire  _wen_T_95 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h2 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_23 = w_valid_s1_0 & _wen_T_95; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5568 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5569 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5570 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5571 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5572 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5573 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5574 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5575 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5576 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5577 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5578 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5579 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5580 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5581 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5582 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5583 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_2_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5584 = 4'h0 == w_addr_s1_0 | _GEN_3440; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5585 = 4'h1 == w_addr_s1_0 | _GEN_3441; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5586 = 4'h2 == w_addr_s1_0 | _GEN_3442; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5587 = 4'h3 == w_addr_s1_0 | _GEN_3443; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5588 = 4'h4 == w_addr_s1_0 | _GEN_3444; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5589 = 4'h5 == w_addr_s1_0 | _GEN_3445; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5590 = 4'h6 == w_addr_s1_0 | _GEN_3446; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5591 = 4'h7 == w_addr_s1_0 | _GEN_3447; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5592 = 4'h8 == w_addr_s1_0 | _GEN_3448; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5593 = 4'h9 == w_addr_s1_0 | _GEN_3449; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5594 = 4'ha == w_addr_s1_0 | _GEN_3450; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5595 = 4'hb == w_addr_s1_0 | _GEN_3451; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5596 = 4'hc == w_addr_s1_0 | _GEN_3452; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5597 = 4'hd == w_addr_s1_0 | _GEN_3453; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5598 = 4'he == w_addr_s1_0 | _GEN_3454; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5599 = 4'hf == w_addr_s1_0 | _GEN_3455; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5600 = wen_23 ? _GEN_5568 : data_0_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5601 = wen_23 ? _GEN_5569 : data_1_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5602 = wen_23 ? _GEN_5570 : data_2_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5603 = wen_23 ? _GEN_5571 : data_3_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5604 = wen_23 ? _GEN_5572 : data_4_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5605 = wen_23 ? _GEN_5573 : data_5_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5606 = wen_23 ? _GEN_5574 : data_6_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5607 = wen_23 ? _GEN_5575 : data_7_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5608 = wen_23 ? _GEN_5576 : data_8_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5609 = wen_23 ? _GEN_5577 : data_9_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5610 = wen_23 ? _GEN_5578 : data_10_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5611 = wen_23 ? _GEN_5579 : data_11_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5612 = wen_23 ? _GEN_5580 : data_12_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5613 = wen_23 ? _GEN_5581 : data_13_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5614 = wen_23 ? _GEN_5582 : data_14_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5615 = wen_23 ? _GEN_5583 : data_15_2_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5616 = wen_23 ? _GEN_5584 : _GEN_3440; // @[Sbuffer.scala 160:18]
  wire  _GEN_5617 = wen_23 ? _GEN_5585 : _GEN_3441; // @[Sbuffer.scala 160:18]
  wire  _GEN_5618 = wen_23 ? _GEN_5586 : _GEN_3442; // @[Sbuffer.scala 160:18]
  wire  _GEN_5619 = wen_23 ? _GEN_5587 : _GEN_3443; // @[Sbuffer.scala 160:18]
  wire  _GEN_5620 = wen_23 ? _GEN_5588 : _GEN_3444; // @[Sbuffer.scala 160:18]
  wire  _GEN_5621 = wen_23 ? _GEN_5589 : _GEN_3445; // @[Sbuffer.scala 160:18]
  wire  _GEN_5622 = wen_23 ? _GEN_5590 : _GEN_3446; // @[Sbuffer.scala 160:18]
  wire  _GEN_5623 = wen_23 ? _GEN_5591 : _GEN_3447; // @[Sbuffer.scala 160:18]
  wire  _GEN_5624 = wen_23 ? _GEN_5592 : _GEN_3448; // @[Sbuffer.scala 160:18]
  wire  _GEN_5625 = wen_23 ? _GEN_5593 : _GEN_3449; // @[Sbuffer.scala 160:18]
  wire  _GEN_5626 = wen_23 ? _GEN_5594 : _GEN_3450; // @[Sbuffer.scala 160:18]
  wire  _GEN_5627 = wen_23 ? _GEN_5595 : _GEN_3451; // @[Sbuffer.scala 160:18]
  wire  _GEN_5628 = wen_23 ? _GEN_5596 : _GEN_3452; // @[Sbuffer.scala 160:18]
  wire  _GEN_5629 = wen_23 ? _GEN_5597 : _GEN_3453; // @[Sbuffer.scala 160:18]
  wire  _GEN_5630 = wen_23 ? _GEN_5598 : _GEN_3454; // @[Sbuffer.scala 160:18]
  wire  _GEN_5631 = wen_23 ? _GEN_5599 : _GEN_3455; // @[Sbuffer.scala 160:18]
  wire  _wen_T_99 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_24 = w_valid_s1_0 & _wen_T_99; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5632 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5633 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5634 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5635 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5636 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5637 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5638 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5639 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5640 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5641 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5642 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5643 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5644 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5645 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5646 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5647 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_3_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5648 = 4'h0 == w_addr_s1_0 | _GEN_3456; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5649 = 4'h1 == w_addr_s1_0 | _GEN_3457; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5650 = 4'h2 == w_addr_s1_0 | _GEN_3458; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5651 = 4'h3 == w_addr_s1_0 | _GEN_3459; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5652 = 4'h4 == w_addr_s1_0 | _GEN_3460; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5653 = 4'h5 == w_addr_s1_0 | _GEN_3461; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5654 = 4'h6 == w_addr_s1_0 | _GEN_3462; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5655 = 4'h7 == w_addr_s1_0 | _GEN_3463; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5656 = 4'h8 == w_addr_s1_0 | _GEN_3464; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5657 = 4'h9 == w_addr_s1_0 | _GEN_3465; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5658 = 4'ha == w_addr_s1_0 | _GEN_3466; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5659 = 4'hb == w_addr_s1_0 | _GEN_3467; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5660 = 4'hc == w_addr_s1_0 | _GEN_3468; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5661 = 4'hd == w_addr_s1_0 | _GEN_3469; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5662 = 4'he == w_addr_s1_0 | _GEN_3470; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5663 = 4'hf == w_addr_s1_0 | _GEN_3471; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5664 = wen_24 ? _GEN_5632 : data_0_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5665 = wen_24 ? _GEN_5633 : data_1_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5666 = wen_24 ? _GEN_5634 : data_2_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5667 = wen_24 ? _GEN_5635 : data_3_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5668 = wen_24 ? _GEN_5636 : data_4_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5669 = wen_24 ? _GEN_5637 : data_5_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5670 = wen_24 ? _GEN_5638 : data_6_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5671 = wen_24 ? _GEN_5639 : data_7_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5672 = wen_24 ? _GEN_5640 : data_8_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5673 = wen_24 ? _GEN_5641 : data_9_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5674 = wen_24 ? _GEN_5642 : data_10_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5675 = wen_24 ? _GEN_5643 : data_11_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5676 = wen_24 ? _GEN_5644 : data_12_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5677 = wen_24 ? _GEN_5645 : data_13_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5678 = wen_24 ? _GEN_5646 : data_14_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5679 = wen_24 ? _GEN_5647 : data_15_3_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5680 = wen_24 ? _GEN_5648 : _GEN_3456; // @[Sbuffer.scala 160:18]
  wire  _GEN_5681 = wen_24 ? _GEN_5649 : _GEN_3457; // @[Sbuffer.scala 160:18]
  wire  _GEN_5682 = wen_24 ? _GEN_5650 : _GEN_3458; // @[Sbuffer.scala 160:18]
  wire  _GEN_5683 = wen_24 ? _GEN_5651 : _GEN_3459; // @[Sbuffer.scala 160:18]
  wire  _GEN_5684 = wen_24 ? _GEN_5652 : _GEN_3460; // @[Sbuffer.scala 160:18]
  wire  _GEN_5685 = wen_24 ? _GEN_5653 : _GEN_3461; // @[Sbuffer.scala 160:18]
  wire  _GEN_5686 = wen_24 ? _GEN_5654 : _GEN_3462; // @[Sbuffer.scala 160:18]
  wire  _GEN_5687 = wen_24 ? _GEN_5655 : _GEN_3463; // @[Sbuffer.scala 160:18]
  wire  _GEN_5688 = wen_24 ? _GEN_5656 : _GEN_3464; // @[Sbuffer.scala 160:18]
  wire  _GEN_5689 = wen_24 ? _GEN_5657 : _GEN_3465; // @[Sbuffer.scala 160:18]
  wire  _GEN_5690 = wen_24 ? _GEN_5658 : _GEN_3466; // @[Sbuffer.scala 160:18]
  wire  _GEN_5691 = wen_24 ? _GEN_5659 : _GEN_3467; // @[Sbuffer.scala 160:18]
  wire  _GEN_5692 = wen_24 ? _GEN_5660 : _GEN_3468; // @[Sbuffer.scala 160:18]
  wire  _GEN_5693 = wen_24 ? _GEN_5661 : _GEN_3469; // @[Sbuffer.scala 160:18]
  wire  _GEN_5694 = wen_24 ? _GEN_5662 : _GEN_3470; // @[Sbuffer.scala 160:18]
  wire  _GEN_5695 = wen_24 ? _GEN_5663 : _GEN_3471; // @[Sbuffer.scala 160:18]
  wire  _wen_T_103 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_25 = w_valid_s1_0 & _wen_T_103; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5696 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5697 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5698 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5699 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5700 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5701 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5702 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5703 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5704 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5705 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5706 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5707 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5708 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5709 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5710 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5711 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_3_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5712 = 4'h0 == w_addr_s1_0 | _GEN_3472; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5713 = 4'h1 == w_addr_s1_0 | _GEN_3473; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5714 = 4'h2 == w_addr_s1_0 | _GEN_3474; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5715 = 4'h3 == w_addr_s1_0 | _GEN_3475; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5716 = 4'h4 == w_addr_s1_0 | _GEN_3476; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5717 = 4'h5 == w_addr_s1_0 | _GEN_3477; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5718 = 4'h6 == w_addr_s1_0 | _GEN_3478; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5719 = 4'h7 == w_addr_s1_0 | _GEN_3479; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5720 = 4'h8 == w_addr_s1_0 | _GEN_3480; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5721 = 4'h9 == w_addr_s1_0 | _GEN_3481; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5722 = 4'ha == w_addr_s1_0 | _GEN_3482; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5723 = 4'hb == w_addr_s1_0 | _GEN_3483; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5724 = 4'hc == w_addr_s1_0 | _GEN_3484; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5725 = 4'hd == w_addr_s1_0 | _GEN_3485; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5726 = 4'he == w_addr_s1_0 | _GEN_3486; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5727 = 4'hf == w_addr_s1_0 | _GEN_3487; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5728 = wen_25 ? _GEN_5696 : data_0_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5729 = wen_25 ? _GEN_5697 : data_1_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5730 = wen_25 ? _GEN_5698 : data_2_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5731 = wen_25 ? _GEN_5699 : data_3_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5732 = wen_25 ? _GEN_5700 : data_4_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5733 = wen_25 ? _GEN_5701 : data_5_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5734 = wen_25 ? _GEN_5702 : data_6_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5735 = wen_25 ? _GEN_5703 : data_7_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5736 = wen_25 ? _GEN_5704 : data_8_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5737 = wen_25 ? _GEN_5705 : data_9_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5738 = wen_25 ? _GEN_5706 : data_10_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5739 = wen_25 ? _GEN_5707 : data_11_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5740 = wen_25 ? _GEN_5708 : data_12_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5741 = wen_25 ? _GEN_5709 : data_13_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5742 = wen_25 ? _GEN_5710 : data_14_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5743 = wen_25 ? _GEN_5711 : data_15_3_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5744 = wen_25 ? _GEN_5712 : _GEN_3472; // @[Sbuffer.scala 160:18]
  wire  _GEN_5745 = wen_25 ? _GEN_5713 : _GEN_3473; // @[Sbuffer.scala 160:18]
  wire  _GEN_5746 = wen_25 ? _GEN_5714 : _GEN_3474; // @[Sbuffer.scala 160:18]
  wire  _GEN_5747 = wen_25 ? _GEN_5715 : _GEN_3475; // @[Sbuffer.scala 160:18]
  wire  _GEN_5748 = wen_25 ? _GEN_5716 : _GEN_3476; // @[Sbuffer.scala 160:18]
  wire  _GEN_5749 = wen_25 ? _GEN_5717 : _GEN_3477; // @[Sbuffer.scala 160:18]
  wire  _GEN_5750 = wen_25 ? _GEN_5718 : _GEN_3478; // @[Sbuffer.scala 160:18]
  wire  _GEN_5751 = wen_25 ? _GEN_5719 : _GEN_3479; // @[Sbuffer.scala 160:18]
  wire  _GEN_5752 = wen_25 ? _GEN_5720 : _GEN_3480; // @[Sbuffer.scala 160:18]
  wire  _GEN_5753 = wen_25 ? _GEN_5721 : _GEN_3481; // @[Sbuffer.scala 160:18]
  wire  _GEN_5754 = wen_25 ? _GEN_5722 : _GEN_3482; // @[Sbuffer.scala 160:18]
  wire  _GEN_5755 = wen_25 ? _GEN_5723 : _GEN_3483; // @[Sbuffer.scala 160:18]
  wire  _GEN_5756 = wen_25 ? _GEN_5724 : _GEN_3484; // @[Sbuffer.scala 160:18]
  wire  _GEN_5757 = wen_25 ? _GEN_5725 : _GEN_3485; // @[Sbuffer.scala 160:18]
  wire  _GEN_5758 = wen_25 ? _GEN_5726 : _GEN_3486; // @[Sbuffer.scala 160:18]
  wire  _GEN_5759 = wen_25 ? _GEN_5727 : _GEN_3487; // @[Sbuffer.scala 160:18]
  wire  _wen_T_107 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_26 = w_valid_s1_0 & _wen_T_107; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5760 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5761 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5762 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5763 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5764 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5765 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5766 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5767 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5768 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5769 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5770 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5771 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5772 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5773 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5774 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5775 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_3_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5776 = 4'h0 == w_addr_s1_0 | _GEN_3488; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5777 = 4'h1 == w_addr_s1_0 | _GEN_3489; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5778 = 4'h2 == w_addr_s1_0 | _GEN_3490; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5779 = 4'h3 == w_addr_s1_0 | _GEN_3491; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5780 = 4'h4 == w_addr_s1_0 | _GEN_3492; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5781 = 4'h5 == w_addr_s1_0 | _GEN_3493; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5782 = 4'h6 == w_addr_s1_0 | _GEN_3494; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5783 = 4'h7 == w_addr_s1_0 | _GEN_3495; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5784 = 4'h8 == w_addr_s1_0 | _GEN_3496; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5785 = 4'h9 == w_addr_s1_0 | _GEN_3497; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5786 = 4'ha == w_addr_s1_0 | _GEN_3498; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5787 = 4'hb == w_addr_s1_0 | _GEN_3499; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5788 = 4'hc == w_addr_s1_0 | _GEN_3500; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5789 = 4'hd == w_addr_s1_0 | _GEN_3501; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5790 = 4'he == w_addr_s1_0 | _GEN_3502; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5791 = 4'hf == w_addr_s1_0 | _GEN_3503; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5792 = wen_26 ? _GEN_5760 : data_0_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5793 = wen_26 ? _GEN_5761 : data_1_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5794 = wen_26 ? _GEN_5762 : data_2_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5795 = wen_26 ? _GEN_5763 : data_3_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5796 = wen_26 ? _GEN_5764 : data_4_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5797 = wen_26 ? _GEN_5765 : data_5_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5798 = wen_26 ? _GEN_5766 : data_6_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5799 = wen_26 ? _GEN_5767 : data_7_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5800 = wen_26 ? _GEN_5768 : data_8_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5801 = wen_26 ? _GEN_5769 : data_9_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5802 = wen_26 ? _GEN_5770 : data_10_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5803 = wen_26 ? _GEN_5771 : data_11_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5804 = wen_26 ? _GEN_5772 : data_12_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5805 = wen_26 ? _GEN_5773 : data_13_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5806 = wen_26 ? _GEN_5774 : data_14_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5807 = wen_26 ? _GEN_5775 : data_15_3_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5808 = wen_26 ? _GEN_5776 : _GEN_3488; // @[Sbuffer.scala 160:18]
  wire  _GEN_5809 = wen_26 ? _GEN_5777 : _GEN_3489; // @[Sbuffer.scala 160:18]
  wire  _GEN_5810 = wen_26 ? _GEN_5778 : _GEN_3490; // @[Sbuffer.scala 160:18]
  wire  _GEN_5811 = wen_26 ? _GEN_5779 : _GEN_3491; // @[Sbuffer.scala 160:18]
  wire  _GEN_5812 = wen_26 ? _GEN_5780 : _GEN_3492; // @[Sbuffer.scala 160:18]
  wire  _GEN_5813 = wen_26 ? _GEN_5781 : _GEN_3493; // @[Sbuffer.scala 160:18]
  wire  _GEN_5814 = wen_26 ? _GEN_5782 : _GEN_3494; // @[Sbuffer.scala 160:18]
  wire  _GEN_5815 = wen_26 ? _GEN_5783 : _GEN_3495; // @[Sbuffer.scala 160:18]
  wire  _GEN_5816 = wen_26 ? _GEN_5784 : _GEN_3496; // @[Sbuffer.scala 160:18]
  wire  _GEN_5817 = wen_26 ? _GEN_5785 : _GEN_3497; // @[Sbuffer.scala 160:18]
  wire  _GEN_5818 = wen_26 ? _GEN_5786 : _GEN_3498; // @[Sbuffer.scala 160:18]
  wire  _GEN_5819 = wen_26 ? _GEN_5787 : _GEN_3499; // @[Sbuffer.scala 160:18]
  wire  _GEN_5820 = wen_26 ? _GEN_5788 : _GEN_3500; // @[Sbuffer.scala 160:18]
  wire  _GEN_5821 = wen_26 ? _GEN_5789 : _GEN_3501; // @[Sbuffer.scala 160:18]
  wire  _GEN_5822 = wen_26 ? _GEN_5790 : _GEN_3502; // @[Sbuffer.scala 160:18]
  wire  _GEN_5823 = wen_26 ? _GEN_5791 : _GEN_3503; // @[Sbuffer.scala 160:18]
  wire  _wen_T_111 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_27 = w_valid_s1_0 & _wen_T_111; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5824 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5825 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5826 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5827 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5828 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5829 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5830 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5831 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5832 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5833 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5834 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5835 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5836 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5837 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5838 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5839 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_3_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5840 = 4'h0 == w_addr_s1_0 | _GEN_3504; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5841 = 4'h1 == w_addr_s1_0 | _GEN_3505; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5842 = 4'h2 == w_addr_s1_0 | _GEN_3506; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5843 = 4'h3 == w_addr_s1_0 | _GEN_3507; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5844 = 4'h4 == w_addr_s1_0 | _GEN_3508; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5845 = 4'h5 == w_addr_s1_0 | _GEN_3509; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5846 = 4'h6 == w_addr_s1_0 | _GEN_3510; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5847 = 4'h7 == w_addr_s1_0 | _GEN_3511; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5848 = 4'h8 == w_addr_s1_0 | _GEN_3512; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5849 = 4'h9 == w_addr_s1_0 | _GEN_3513; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5850 = 4'ha == w_addr_s1_0 | _GEN_3514; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5851 = 4'hb == w_addr_s1_0 | _GEN_3515; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5852 = 4'hc == w_addr_s1_0 | _GEN_3516; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5853 = 4'hd == w_addr_s1_0 | _GEN_3517; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5854 = 4'he == w_addr_s1_0 | _GEN_3518; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5855 = 4'hf == w_addr_s1_0 | _GEN_3519; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5856 = wen_27 ? _GEN_5824 : data_0_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5857 = wen_27 ? _GEN_5825 : data_1_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5858 = wen_27 ? _GEN_5826 : data_2_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5859 = wen_27 ? _GEN_5827 : data_3_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5860 = wen_27 ? _GEN_5828 : data_4_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5861 = wen_27 ? _GEN_5829 : data_5_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5862 = wen_27 ? _GEN_5830 : data_6_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5863 = wen_27 ? _GEN_5831 : data_7_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5864 = wen_27 ? _GEN_5832 : data_8_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5865 = wen_27 ? _GEN_5833 : data_9_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5866 = wen_27 ? _GEN_5834 : data_10_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5867 = wen_27 ? _GEN_5835 : data_11_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5868 = wen_27 ? _GEN_5836 : data_12_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5869 = wen_27 ? _GEN_5837 : data_13_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5870 = wen_27 ? _GEN_5838 : data_14_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5871 = wen_27 ? _GEN_5839 : data_15_3_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5872 = wen_27 ? _GEN_5840 : _GEN_3504; // @[Sbuffer.scala 160:18]
  wire  _GEN_5873 = wen_27 ? _GEN_5841 : _GEN_3505; // @[Sbuffer.scala 160:18]
  wire  _GEN_5874 = wen_27 ? _GEN_5842 : _GEN_3506; // @[Sbuffer.scala 160:18]
  wire  _GEN_5875 = wen_27 ? _GEN_5843 : _GEN_3507; // @[Sbuffer.scala 160:18]
  wire  _GEN_5876 = wen_27 ? _GEN_5844 : _GEN_3508; // @[Sbuffer.scala 160:18]
  wire  _GEN_5877 = wen_27 ? _GEN_5845 : _GEN_3509; // @[Sbuffer.scala 160:18]
  wire  _GEN_5878 = wen_27 ? _GEN_5846 : _GEN_3510; // @[Sbuffer.scala 160:18]
  wire  _GEN_5879 = wen_27 ? _GEN_5847 : _GEN_3511; // @[Sbuffer.scala 160:18]
  wire  _GEN_5880 = wen_27 ? _GEN_5848 : _GEN_3512; // @[Sbuffer.scala 160:18]
  wire  _GEN_5881 = wen_27 ? _GEN_5849 : _GEN_3513; // @[Sbuffer.scala 160:18]
  wire  _GEN_5882 = wen_27 ? _GEN_5850 : _GEN_3514; // @[Sbuffer.scala 160:18]
  wire  _GEN_5883 = wen_27 ? _GEN_5851 : _GEN_3515; // @[Sbuffer.scala 160:18]
  wire  _GEN_5884 = wen_27 ? _GEN_5852 : _GEN_3516; // @[Sbuffer.scala 160:18]
  wire  _GEN_5885 = wen_27 ? _GEN_5853 : _GEN_3517; // @[Sbuffer.scala 160:18]
  wire  _GEN_5886 = wen_27 ? _GEN_5854 : _GEN_3518; // @[Sbuffer.scala 160:18]
  wire  _GEN_5887 = wen_27 ? _GEN_5855 : _GEN_3519; // @[Sbuffer.scala 160:18]
  wire  _wen_T_115 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_28 = w_valid_s1_0 & _wen_T_115; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5888 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5889 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5890 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5891 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5892 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5893 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5894 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5895 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5896 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5897 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5898 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5899 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5900 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5901 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5902 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5903 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_3_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5904 = 4'h0 == w_addr_s1_0 | _GEN_3520; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5905 = 4'h1 == w_addr_s1_0 | _GEN_3521; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5906 = 4'h2 == w_addr_s1_0 | _GEN_3522; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5907 = 4'h3 == w_addr_s1_0 | _GEN_3523; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5908 = 4'h4 == w_addr_s1_0 | _GEN_3524; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5909 = 4'h5 == w_addr_s1_0 | _GEN_3525; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5910 = 4'h6 == w_addr_s1_0 | _GEN_3526; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5911 = 4'h7 == w_addr_s1_0 | _GEN_3527; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5912 = 4'h8 == w_addr_s1_0 | _GEN_3528; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5913 = 4'h9 == w_addr_s1_0 | _GEN_3529; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5914 = 4'ha == w_addr_s1_0 | _GEN_3530; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5915 = 4'hb == w_addr_s1_0 | _GEN_3531; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5916 = 4'hc == w_addr_s1_0 | _GEN_3532; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5917 = 4'hd == w_addr_s1_0 | _GEN_3533; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5918 = 4'he == w_addr_s1_0 | _GEN_3534; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5919 = 4'hf == w_addr_s1_0 | _GEN_3535; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5920 = wen_28 ? _GEN_5888 : data_0_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5921 = wen_28 ? _GEN_5889 : data_1_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5922 = wen_28 ? _GEN_5890 : data_2_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5923 = wen_28 ? _GEN_5891 : data_3_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5924 = wen_28 ? _GEN_5892 : data_4_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5925 = wen_28 ? _GEN_5893 : data_5_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5926 = wen_28 ? _GEN_5894 : data_6_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5927 = wen_28 ? _GEN_5895 : data_7_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5928 = wen_28 ? _GEN_5896 : data_8_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5929 = wen_28 ? _GEN_5897 : data_9_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5930 = wen_28 ? _GEN_5898 : data_10_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5931 = wen_28 ? _GEN_5899 : data_11_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5932 = wen_28 ? _GEN_5900 : data_12_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5933 = wen_28 ? _GEN_5901 : data_13_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5934 = wen_28 ? _GEN_5902 : data_14_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5935 = wen_28 ? _GEN_5903 : data_15_3_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_5936 = wen_28 ? _GEN_5904 : _GEN_3520; // @[Sbuffer.scala 160:18]
  wire  _GEN_5937 = wen_28 ? _GEN_5905 : _GEN_3521; // @[Sbuffer.scala 160:18]
  wire  _GEN_5938 = wen_28 ? _GEN_5906 : _GEN_3522; // @[Sbuffer.scala 160:18]
  wire  _GEN_5939 = wen_28 ? _GEN_5907 : _GEN_3523; // @[Sbuffer.scala 160:18]
  wire  _GEN_5940 = wen_28 ? _GEN_5908 : _GEN_3524; // @[Sbuffer.scala 160:18]
  wire  _GEN_5941 = wen_28 ? _GEN_5909 : _GEN_3525; // @[Sbuffer.scala 160:18]
  wire  _GEN_5942 = wen_28 ? _GEN_5910 : _GEN_3526; // @[Sbuffer.scala 160:18]
  wire  _GEN_5943 = wen_28 ? _GEN_5911 : _GEN_3527; // @[Sbuffer.scala 160:18]
  wire  _GEN_5944 = wen_28 ? _GEN_5912 : _GEN_3528; // @[Sbuffer.scala 160:18]
  wire  _GEN_5945 = wen_28 ? _GEN_5913 : _GEN_3529; // @[Sbuffer.scala 160:18]
  wire  _GEN_5946 = wen_28 ? _GEN_5914 : _GEN_3530; // @[Sbuffer.scala 160:18]
  wire  _GEN_5947 = wen_28 ? _GEN_5915 : _GEN_3531; // @[Sbuffer.scala 160:18]
  wire  _GEN_5948 = wen_28 ? _GEN_5916 : _GEN_3532; // @[Sbuffer.scala 160:18]
  wire  _GEN_5949 = wen_28 ? _GEN_5917 : _GEN_3533; // @[Sbuffer.scala 160:18]
  wire  _GEN_5950 = wen_28 ? _GEN_5918 : _GEN_3534; // @[Sbuffer.scala 160:18]
  wire  _GEN_5951 = wen_28 ? _GEN_5919 : _GEN_3535; // @[Sbuffer.scala 160:18]
  wire  _wen_T_119 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_29 = w_valid_s1_0 & _wen_T_119; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_5952 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5953 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5954 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5955 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5956 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5957 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5958 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5959 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5960 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5961 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5962 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5963 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5964 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5965 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5966 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_5967 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_3_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_5968 = 4'h0 == w_addr_s1_0 | _GEN_3536; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5969 = 4'h1 == w_addr_s1_0 | _GEN_3537; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5970 = 4'h2 == w_addr_s1_0 | _GEN_3538; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5971 = 4'h3 == w_addr_s1_0 | _GEN_3539; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5972 = 4'h4 == w_addr_s1_0 | _GEN_3540; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5973 = 4'h5 == w_addr_s1_0 | _GEN_3541; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5974 = 4'h6 == w_addr_s1_0 | _GEN_3542; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5975 = 4'h7 == w_addr_s1_0 | _GEN_3543; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5976 = 4'h8 == w_addr_s1_0 | _GEN_3544; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5977 = 4'h9 == w_addr_s1_0 | _GEN_3545; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5978 = 4'ha == w_addr_s1_0 | _GEN_3546; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5979 = 4'hb == w_addr_s1_0 | _GEN_3547; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5980 = 4'hc == w_addr_s1_0 | _GEN_3548; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5981 = 4'hd == w_addr_s1_0 | _GEN_3549; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5982 = 4'he == w_addr_s1_0 | _GEN_3550; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_5983 = 4'hf == w_addr_s1_0 | _GEN_3551; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_5984 = wen_29 ? _GEN_5952 : data_0_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5985 = wen_29 ? _GEN_5953 : data_1_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5986 = wen_29 ? _GEN_5954 : data_2_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5987 = wen_29 ? _GEN_5955 : data_3_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5988 = wen_29 ? _GEN_5956 : data_4_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5989 = wen_29 ? _GEN_5957 : data_5_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5990 = wen_29 ? _GEN_5958 : data_6_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5991 = wen_29 ? _GEN_5959 : data_7_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5992 = wen_29 ? _GEN_5960 : data_8_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5993 = wen_29 ? _GEN_5961 : data_9_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5994 = wen_29 ? _GEN_5962 : data_10_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5995 = wen_29 ? _GEN_5963 : data_11_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5996 = wen_29 ? _GEN_5964 : data_12_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5997 = wen_29 ? _GEN_5965 : data_13_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5998 = wen_29 ? _GEN_5966 : data_14_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_5999 = wen_29 ? _GEN_5967 : data_15_3_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6000 = wen_29 ? _GEN_5968 : _GEN_3536; // @[Sbuffer.scala 160:18]
  wire  _GEN_6001 = wen_29 ? _GEN_5969 : _GEN_3537; // @[Sbuffer.scala 160:18]
  wire  _GEN_6002 = wen_29 ? _GEN_5970 : _GEN_3538; // @[Sbuffer.scala 160:18]
  wire  _GEN_6003 = wen_29 ? _GEN_5971 : _GEN_3539; // @[Sbuffer.scala 160:18]
  wire  _GEN_6004 = wen_29 ? _GEN_5972 : _GEN_3540; // @[Sbuffer.scala 160:18]
  wire  _GEN_6005 = wen_29 ? _GEN_5973 : _GEN_3541; // @[Sbuffer.scala 160:18]
  wire  _GEN_6006 = wen_29 ? _GEN_5974 : _GEN_3542; // @[Sbuffer.scala 160:18]
  wire  _GEN_6007 = wen_29 ? _GEN_5975 : _GEN_3543; // @[Sbuffer.scala 160:18]
  wire  _GEN_6008 = wen_29 ? _GEN_5976 : _GEN_3544; // @[Sbuffer.scala 160:18]
  wire  _GEN_6009 = wen_29 ? _GEN_5977 : _GEN_3545; // @[Sbuffer.scala 160:18]
  wire  _GEN_6010 = wen_29 ? _GEN_5978 : _GEN_3546; // @[Sbuffer.scala 160:18]
  wire  _GEN_6011 = wen_29 ? _GEN_5979 : _GEN_3547; // @[Sbuffer.scala 160:18]
  wire  _GEN_6012 = wen_29 ? _GEN_5980 : _GEN_3548; // @[Sbuffer.scala 160:18]
  wire  _GEN_6013 = wen_29 ? _GEN_5981 : _GEN_3549; // @[Sbuffer.scala 160:18]
  wire  _GEN_6014 = wen_29 ? _GEN_5982 : _GEN_3550; // @[Sbuffer.scala 160:18]
  wire  _GEN_6015 = wen_29 ? _GEN_5983 : _GEN_3551; // @[Sbuffer.scala 160:18]
  wire  _wen_T_123 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_30 = w_valid_s1_0 & _wen_T_123; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6016 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6017 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6018 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6019 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6020 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6021 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6022 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6023 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6024 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6025 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6026 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6027 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6028 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6029 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6030 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6031 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_3_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6032 = 4'h0 == w_addr_s1_0 | _GEN_3552; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6033 = 4'h1 == w_addr_s1_0 | _GEN_3553; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6034 = 4'h2 == w_addr_s1_0 | _GEN_3554; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6035 = 4'h3 == w_addr_s1_0 | _GEN_3555; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6036 = 4'h4 == w_addr_s1_0 | _GEN_3556; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6037 = 4'h5 == w_addr_s1_0 | _GEN_3557; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6038 = 4'h6 == w_addr_s1_0 | _GEN_3558; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6039 = 4'h7 == w_addr_s1_0 | _GEN_3559; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6040 = 4'h8 == w_addr_s1_0 | _GEN_3560; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6041 = 4'h9 == w_addr_s1_0 | _GEN_3561; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6042 = 4'ha == w_addr_s1_0 | _GEN_3562; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6043 = 4'hb == w_addr_s1_0 | _GEN_3563; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6044 = 4'hc == w_addr_s1_0 | _GEN_3564; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6045 = 4'hd == w_addr_s1_0 | _GEN_3565; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6046 = 4'he == w_addr_s1_0 | _GEN_3566; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6047 = 4'hf == w_addr_s1_0 | _GEN_3567; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6048 = wen_30 ? _GEN_6016 : data_0_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6049 = wen_30 ? _GEN_6017 : data_1_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6050 = wen_30 ? _GEN_6018 : data_2_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6051 = wen_30 ? _GEN_6019 : data_3_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6052 = wen_30 ? _GEN_6020 : data_4_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6053 = wen_30 ? _GEN_6021 : data_5_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6054 = wen_30 ? _GEN_6022 : data_6_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6055 = wen_30 ? _GEN_6023 : data_7_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6056 = wen_30 ? _GEN_6024 : data_8_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6057 = wen_30 ? _GEN_6025 : data_9_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6058 = wen_30 ? _GEN_6026 : data_10_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6059 = wen_30 ? _GEN_6027 : data_11_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6060 = wen_30 ? _GEN_6028 : data_12_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6061 = wen_30 ? _GEN_6029 : data_13_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6062 = wen_30 ? _GEN_6030 : data_14_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6063 = wen_30 ? _GEN_6031 : data_15_3_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6064 = wen_30 ? _GEN_6032 : _GEN_3552; // @[Sbuffer.scala 160:18]
  wire  _GEN_6065 = wen_30 ? _GEN_6033 : _GEN_3553; // @[Sbuffer.scala 160:18]
  wire  _GEN_6066 = wen_30 ? _GEN_6034 : _GEN_3554; // @[Sbuffer.scala 160:18]
  wire  _GEN_6067 = wen_30 ? _GEN_6035 : _GEN_3555; // @[Sbuffer.scala 160:18]
  wire  _GEN_6068 = wen_30 ? _GEN_6036 : _GEN_3556; // @[Sbuffer.scala 160:18]
  wire  _GEN_6069 = wen_30 ? _GEN_6037 : _GEN_3557; // @[Sbuffer.scala 160:18]
  wire  _GEN_6070 = wen_30 ? _GEN_6038 : _GEN_3558; // @[Sbuffer.scala 160:18]
  wire  _GEN_6071 = wen_30 ? _GEN_6039 : _GEN_3559; // @[Sbuffer.scala 160:18]
  wire  _GEN_6072 = wen_30 ? _GEN_6040 : _GEN_3560; // @[Sbuffer.scala 160:18]
  wire  _GEN_6073 = wen_30 ? _GEN_6041 : _GEN_3561; // @[Sbuffer.scala 160:18]
  wire  _GEN_6074 = wen_30 ? _GEN_6042 : _GEN_3562; // @[Sbuffer.scala 160:18]
  wire  _GEN_6075 = wen_30 ? _GEN_6043 : _GEN_3563; // @[Sbuffer.scala 160:18]
  wire  _GEN_6076 = wen_30 ? _GEN_6044 : _GEN_3564; // @[Sbuffer.scala 160:18]
  wire  _GEN_6077 = wen_30 ? _GEN_6045 : _GEN_3565; // @[Sbuffer.scala 160:18]
  wire  _GEN_6078 = wen_30 ? _GEN_6046 : _GEN_3566; // @[Sbuffer.scala 160:18]
  wire  _GEN_6079 = wen_30 ? _GEN_6047 : _GEN_3567; // @[Sbuffer.scala 160:18]
  wire  _wen_T_127 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h3 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_31 = w_valid_s1_0 & _wen_T_127; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6080 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6081 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6082 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6083 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6084 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6085 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6086 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6087 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6088 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6089 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6090 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6091 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6092 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6093 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6094 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6095 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_3_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6096 = 4'h0 == w_addr_s1_0 | _GEN_3568; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6097 = 4'h1 == w_addr_s1_0 | _GEN_3569; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6098 = 4'h2 == w_addr_s1_0 | _GEN_3570; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6099 = 4'h3 == w_addr_s1_0 | _GEN_3571; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6100 = 4'h4 == w_addr_s1_0 | _GEN_3572; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6101 = 4'h5 == w_addr_s1_0 | _GEN_3573; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6102 = 4'h6 == w_addr_s1_0 | _GEN_3574; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6103 = 4'h7 == w_addr_s1_0 | _GEN_3575; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6104 = 4'h8 == w_addr_s1_0 | _GEN_3576; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6105 = 4'h9 == w_addr_s1_0 | _GEN_3577; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6106 = 4'ha == w_addr_s1_0 | _GEN_3578; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6107 = 4'hb == w_addr_s1_0 | _GEN_3579; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6108 = 4'hc == w_addr_s1_0 | _GEN_3580; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6109 = 4'hd == w_addr_s1_0 | _GEN_3581; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6110 = 4'he == w_addr_s1_0 | _GEN_3582; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6111 = 4'hf == w_addr_s1_0 | _GEN_3583; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6112 = wen_31 ? _GEN_6080 : data_0_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6113 = wen_31 ? _GEN_6081 : data_1_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6114 = wen_31 ? _GEN_6082 : data_2_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6115 = wen_31 ? _GEN_6083 : data_3_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6116 = wen_31 ? _GEN_6084 : data_4_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6117 = wen_31 ? _GEN_6085 : data_5_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6118 = wen_31 ? _GEN_6086 : data_6_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6119 = wen_31 ? _GEN_6087 : data_7_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6120 = wen_31 ? _GEN_6088 : data_8_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6121 = wen_31 ? _GEN_6089 : data_9_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6122 = wen_31 ? _GEN_6090 : data_10_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6123 = wen_31 ? _GEN_6091 : data_11_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6124 = wen_31 ? _GEN_6092 : data_12_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6125 = wen_31 ? _GEN_6093 : data_13_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6126 = wen_31 ? _GEN_6094 : data_14_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6127 = wen_31 ? _GEN_6095 : data_15_3_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6128 = wen_31 ? _GEN_6096 : _GEN_3568; // @[Sbuffer.scala 160:18]
  wire  _GEN_6129 = wen_31 ? _GEN_6097 : _GEN_3569; // @[Sbuffer.scala 160:18]
  wire  _GEN_6130 = wen_31 ? _GEN_6098 : _GEN_3570; // @[Sbuffer.scala 160:18]
  wire  _GEN_6131 = wen_31 ? _GEN_6099 : _GEN_3571; // @[Sbuffer.scala 160:18]
  wire  _GEN_6132 = wen_31 ? _GEN_6100 : _GEN_3572; // @[Sbuffer.scala 160:18]
  wire  _GEN_6133 = wen_31 ? _GEN_6101 : _GEN_3573; // @[Sbuffer.scala 160:18]
  wire  _GEN_6134 = wen_31 ? _GEN_6102 : _GEN_3574; // @[Sbuffer.scala 160:18]
  wire  _GEN_6135 = wen_31 ? _GEN_6103 : _GEN_3575; // @[Sbuffer.scala 160:18]
  wire  _GEN_6136 = wen_31 ? _GEN_6104 : _GEN_3576; // @[Sbuffer.scala 160:18]
  wire  _GEN_6137 = wen_31 ? _GEN_6105 : _GEN_3577; // @[Sbuffer.scala 160:18]
  wire  _GEN_6138 = wen_31 ? _GEN_6106 : _GEN_3578; // @[Sbuffer.scala 160:18]
  wire  _GEN_6139 = wen_31 ? _GEN_6107 : _GEN_3579; // @[Sbuffer.scala 160:18]
  wire  _GEN_6140 = wen_31 ? _GEN_6108 : _GEN_3580; // @[Sbuffer.scala 160:18]
  wire  _GEN_6141 = wen_31 ? _GEN_6109 : _GEN_3581; // @[Sbuffer.scala 160:18]
  wire  _GEN_6142 = wen_31 ? _GEN_6110 : _GEN_3582; // @[Sbuffer.scala 160:18]
  wire  _GEN_6143 = wen_31 ? _GEN_6111 : _GEN_3583; // @[Sbuffer.scala 160:18]
  wire  _wen_T_131 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_32 = w_valid_s1_0 & _wen_T_131; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6144 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6145 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6146 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6147 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6148 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6149 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6150 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6151 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6152 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6153 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6154 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6155 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6156 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6157 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6158 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6159 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_4_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6160 = 4'h0 == w_addr_s1_0 | _GEN_3584; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6161 = 4'h1 == w_addr_s1_0 | _GEN_3585; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6162 = 4'h2 == w_addr_s1_0 | _GEN_3586; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6163 = 4'h3 == w_addr_s1_0 | _GEN_3587; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6164 = 4'h4 == w_addr_s1_0 | _GEN_3588; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6165 = 4'h5 == w_addr_s1_0 | _GEN_3589; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6166 = 4'h6 == w_addr_s1_0 | _GEN_3590; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6167 = 4'h7 == w_addr_s1_0 | _GEN_3591; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6168 = 4'h8 == w_addr_s1_0 | _GEN_3592; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6169 = 4'h9 == w_addr_s1_0 | _GEN_3593; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6170 = 4'ha == w_addr_s1_0 | _GEN_3594; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6171 = 4'hb == w_addr_s1_0 | _GEN_3595; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6172 = 4'hc == w_addr_s1_0 | _GEN_3596; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6173 = 4'hd == w_addr_s1_0 | _GEN_3597; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6174 = 4'he == w_addr_s1_0 | _GEN_3598; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6175 = 4'hf == w_addr_s1_0 | _GEN_3599; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6176 = wen_32 ? _GEN_6144 : data_0_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6177 = wen_32 ? _GEN_6145 : data_1_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6178 = wen_32 ? _GEN_6146 : data_2_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6179 = wen_32 ? _GEN_6147 : data_3_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6180 = wen_32 ? _GEN_6148 : data_4_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6181 = wen_32 ? _GEN_6149 : data_5_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6182 = wen_32 ? _GEN_6150 : data_6_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6183 = wen_32 ? _GEN_6151 : data_7_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6184 = wen_32 ? _GEN_6152 : data_8_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6185 = wen_32 ? _GEN_6153 : data_9_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6186 = wen_32 ? _GEN_6154 : data_10_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6187 = wen_32 ? _GEN_6155 : data_11_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6188 = wen_32 ? _GEN_6156 : data_12_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6189 = wen_32 ? _GEN_6157 : data_13_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6190 = wen_32 ? _GEN_6158 : data_14_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6191 = wen_32 ? _GEN_6159 : data_15_4_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6192 = wen_32 ? _GEN_6160 : _GEN_3584; // @[Sbuffer.scala 160:18]
  wire  _GEN_6193 = wen_32 ? _GEN_6161 : _GEN_3585; // @[Sbuffer.scala 160:18]
  wire  _GEN_6194 = wen_32 ? _GEN_6162 : _GEN_3586; // @[Sbuffer.scala 160:18]
  wire  _GEN_6195 = wen_32 ? _GEN_6163 : _GEN_3587; // @[Sbuffer.scala 160:18]
  wire  _GEN_6196 = wen_32 ? _GEN_6164 : _GEN_3588; // @[Sbuffer.scala 160:18]
  wire  _GEN_6197 = wen_32 ? _GEN_6165 : _GEN_3589; // @[Sbuffer.scala 160:18]
  wire  _GEN_6198 = wen_32 ? _GEN_6166 : _GEN_3590; // @[Sbuffer.scala 160:18]
  wire  _GEN_6199 = wen_32 ? _GEN_6167 : _GEN_3591; // @[Sbuffer.scala 160:18]
  wire  _GEN_6200 = wen_32 ? _GEN_6168 : _GEN_3592; // @[Sbuffer.scala 160:18]
  wire  _GEN_6201 = wen_32 ? _GEN_6169 : _GEN_3593; // @[Sbuffer.scala 160:18]
  wire  _GEN_6202 = wen_32 ? _GEN_6170 : _GEN_3594; // @[Sbuffer.scala 160:18]
  wire  _GEN_6203 = wen_32 ? _GEN_6171 : _GEN_3595; // @[Sbuffer.scala 160:18]
  wire  _GEN_6204 = wen_32 ? _GEN_6172 : _GEN_3596; // @[Sbuffer.scala 160:18]
  wire  _GEN_6205 = wen_32 ? _GEN_6173 : _GEN_3597; // @[Sbuffer.scala 160:18]
  wire  _GEN_6206 = wen_32 ? _GEN_6174 : _GEN_3598; // @[Sbuffer.scala 160:18]
  wire  _GEN_6207 = wen_32 ? _GEN_6175 : _GEN_3599; // @[Sbuffer.scala 160:18]
  wire  _wen_T_135 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_33 = w_valid_s1_0 & _wen_T_135; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6208 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6209 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6210 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6211 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6212 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6213 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6214 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6215 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6216 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6217 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6218 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6219 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6220 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6221 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6222 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6223 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_4_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6224 = 4'h0 == w_addr_s1_0 | _GEN_3600; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6225 = 4'h1 == w_addr_s1_0 | _GEN_3601; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6226 = 4'h2 == w_addr_s1_0 | _GEN_3602; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6227 = 4'h3 == w_addr_s1_0 | _GEN_3603; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6228 = 4'h4 == w_addr_s1_0 | _GEN_3604; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6229 = 4'h5 == w_addr_s1_0 | _GEN_3605; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6230 = 4'h6 == w_addr_s1_0 | _GEN_3606; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6231 = 4'h7 == w_addr_s1_0 | _GEN_3607; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6232 = 4'h8 == w_addr_s1_0 | _GEN_3608; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6233 = 4'h9 == w_addr_s1_0 | _GEN_3609; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6234 = 4'ha == w_addr_s1_0 | _GEN_3610; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6235 = 4'hb == w_addr_s1_0 | _GEN_3611; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6236 = 4'hc == w_addr_s1_0 | _GEN_3612; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6237 = 4'hd == w_addr_s1_0 | _GEN_3613; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6238 = 4'he == w_addr_s1_0 | _GEN_3614; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6239 = 4'hf == w_addr_s1_0 | _GEN_3615; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6240 = wen_33 ? _GEN_6208 : data_0_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6241 = wen_33 ? _GEN_6209 : data_1_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6242 = wen_33 ? _GEN_6210 : data_2_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6243 = wen_33 ? _GEN_6211 : data_3_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6244 = wen_33 ? _GEN_6212 : data_4_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6245 = wen_33 ? _GEN_6213 : data_5_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6246 = wen_33 ? _GEN_6214 : data_6_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6247 = wen_33 ? _GEN_6215 : data_7_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6248 = wen_33 ? _GEN_6216 : data_8_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6249 = wen_33 ? _GEN_6217 : data_9_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6250 = wen_33 ? _GEN_6218 : data_10_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6251 = wen_33 ? _GEN_6219 : data_11_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6252 = wen_33 ? _GEN_6220 : data_12_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6253 = wen_33 ? _GEN_6221 : data_13_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6254 = wen_33 ? _GEN_6222 : data_14_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6255 = wen_33 ? _GEN_6223 : data_15_4_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6256 = wen_33 ? _GEN_6224 : _GEN_3600; // @[Sbuffer.scala 160:18]
  wire  _GEN_6257 = wen_33 ? _GEN_6225 : _GEN_3601; // @[Sbuffer.scala 160:18]
  wire  _GEN_6258 = wen_33 ? _GEN_6226 : _GEN_3602; // @[Sbuffer.scala 160:18]
  wire  _GEN_6259 = wen_33 ? _GEN_6227 : _GEN_3603; // @[Sbuffer.scala 160:18]
  wire  _GEN_6260 = wen_33 ? _GEN_6228 : _GEN_3604; // @[Sbuffer.scala 160:18]
  wire  _GEN_6261 = wen_33 ? _GEN_6229 : _GEN_3605; // @[Sbuffer.scala 160:18]
  wire  _GEN_6262 = wen_33 ? _GEN_6230 : _GEN_3606; // @[Sbuffer.scala 160:18]
  wire  _GEN_6263 = wen_33 ? _GEN_6231 : _GEN_3607; // @[Sbuffer.scala 160:18]
  wire  _GEN_6264 = wen_33 ? _GEN_6232 : _GEN_3608; // @[Sbuffer.scala 160:18]
  wire  _GEN_6265 = wen_33 ? _GEN_6233 : _GEN_3609; // @[Sbuffer.scala 160:18]
  wire  _GEN_6266 = wen_33 ? _GEN_6234 : _GEN_3610; // @[Sbuffer.scala 160:18]
  wire  _GEN_6267 = wen_33 ? _GEN_6235 : _GEN_3611; // @[Sbuffer.scala 160:18]
  wire  _GEN_6268 = wen_33 ? _GEN_6236 : _GEN_3612; // @[Sbuffer.scala 160:18]
  wire  _GEN_6269 = wen_33 ? _GEN_6237 : _GEN_3613; // @[Sbuffer.scala 160:18]
  wire  _GEN_6270 = wen_33 ? _GEN_6238 : _GEN_3614; // @[Sbuffer.scala 160:18]
  wire  _GEN_6271 = wen_33 ? _GEN_6239 : _GEN_3615; // @[Sbuffer.scala 160:18]
  wire  _wen_T_139 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_34 = w_valid_s1_0 & _wen_T_139; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6272 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6273 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6274 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6275 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6276 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6277 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6278 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6279 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6280 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6281 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6282 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6283 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6284 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6285 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6286 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6287 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_4_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6288 = 4'h0 == w_addr_s1_0 | _GEN_3616; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6289 = 4'h1 == w_addr_s1_0 | _GEN_3617; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6290 = 4'h2 == w_addr_s1_0 | _GEN_3618; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6291 = 4'h3 == w_addr_s1_0 | _GEN_3619; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6292 = 4'h4 == w_addr_s1_0 | _GEN_3620; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6293 = 4'h5 == w_addr_s1_0 | _GEN_3621; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6294 = 4'h6 == w_addr_s1_0 | _GEN_3622; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6295 = 4'h7 == w_addr_s1_0 | _GEN_3623; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6296 = 4'h8 == w_addr_s1_0 | _GEN_3624; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6297 = 4'h9 == w_addr_s1_0 | _GEN_3625; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6298 = 4'ha == w_addr_s1_0 | _GEN_3626; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6299 = 4'hb == w_addr_s1_0 | _GEN_3627; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6300 = 4'hc == w_addr_s1_0 | _GEN_3628; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6301 = 4'hd == w_addr_s1_0 | _GEN_3629; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6302 = 4'he == w_addr_s1_0 | _GEN_3630; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6303 = 4'hf == w_addr_s1_0 | _GEN_3631; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6304 = wen_34 ? _GEN_6272 : data_0_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6305 = wen_34 ? _GEN_6273 : data_1_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6306 = wen_34 ? _GEN_6274 : data_2_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6307 = wen_34 ? _GEN_6275 : data_3_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6308 = wen_34 ? _GEN_6276 : data_4_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6309 = wen_34 ? _GEN_6277 : data_5_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6310 = wen_34 ? _GEN_6278 : data_6_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6311 = wen_34 ? _GEN_6279 : data_7_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6312 = wen_34 ? _GEN_6280 : data_8_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6313 = wen_34 ? _GEN_6281 : data_9_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6314 = wen_34 ? _GEN_6282 : data_10_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6315 = wen_34 ? _GEN_6283 : data_11_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6316 = wen_34 ? _GEN_6284 : data_12_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6317 = wen_34 ? _GEN_6285 : data_13_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6318 = wen_34 ? _GEN_6286 : data_14_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6319 = wen_34 ? _GEN_6287 : data_15_4_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6320 = wen_34 ? _GEN_6288 : _GEN_3616; // @[Sbuffer.scala 160:18]
  wire  _GEN_6321 = wen_34 ? _GEN_6289 : _GEN_3617; // @[Sbuffer.scala 160:18]
  wire  _GEN_6322 = wen_34 ? _GEN_6290 : _GEN_3618; // @[Sbuffer.scala 160:18]
  wire  _GEN_6323 = wen_34 ? _GEN_6291 : _GEN_3619; // @[Sbuffer.scala 160:18]
  wire  _GEN_6324 = wen_34 ? _GEN_6292 : _GEN_3620; // @[Sbuffer.scala 160:18]
  wire  _GEN_6325 = wen_34 ? _GEN_6293 : _GEN_3621; // @[Sbuffer.scala 160:18]
  wire  _GEN_6326 = wen_34 ? _GEN_6294 : _GEN_3622; // @[Sbuffer.scala 160:18]
  wire  _GEN_6327 = wen_34 ? _GEN_6295 : _GEN_3623; // @[Sbuffer.scala 160:18]
  wire  _GEN_6328 = wen_34 ? _GEN_6296 : _GEN_3624; // @[Sbuffer.scala 160:18]
  wire  _GEN_6329 = wen_34 ? _GEN_6297 : _GEN_3625; // @[Sbuffer.scala 160:18]
  wire  _GEN_6330 = wen_34 ? _GEN_6298 : _GEN_3626; // @[Sbuffer.scala 160:18]
  wire  _GEN_6331 = wen_34 ? _GEN_6299 : _GEN_3627; // @[Sbuffer.scala 160:18]
  wire  _GEN_6332 = wen_34 ? _GEN_6300 : _GEN_3628; // @[Sbuffer.scala 160:18]
  wire  _GEN_6333 = wen_34 ? _GEN_6301 : _GEN_3629; // @[Sbuffer.scala 160:18]
  wire  _GEN_6334 = wen_34 ? _GEN_6302 : _GEN_3630; // @[Sbuffer.scala 160:18]
  wire  _GEN_6335 = wen_34 ? _GEN_6303 : _GEN_3631; // @[Sbuffer.scala 160:18]
  wire  _wen_T_143 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_35 = w_valid_s1_0 & _wen_T_143; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6336 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6337 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6338 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6339 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6340 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6341 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6342 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6343 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6344 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6345 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6346 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6347 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6348 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6349 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6350 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6351 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_4_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6352 = 4'h0 == w_addr_s1_0 | _GEN_3632; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6353 = 4'h1 == w_addr_s1_0 | _GEN_3633; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6354 = 4'h2 == w_addr_s1_0 | _GEN_3634; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6355 = 4'h3 == w_addr_s1_0 | _GEN_3635; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6356 = 4'h4 == w_addr_s1_0 | _GEN_3636; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6357 = 4'h5 == w_addr_s1_0 | _GEN_3637; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6358 = 4'h6 == w_addr_s1_0 | _GEN_3638; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6359 = 4'h7 == w_addr_s1_0 | _GEN_3639; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6360 = 4'h8 == w_addr_s1_0 | _GEN_3640; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6361 = 4'h9 == w_addr_s1_0 | _GEN_3641; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6362 = 4'ha == w_addr_s1_0 | _GEN_3642; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6363 = 4'hb == w_addr_s1_0 | _GEN_3643; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6364 = 4'hc == w_addr_s1_0 | _GEN_3644; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6365 = 4'hd == w_addr_s1_0 | _GEN_3645; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6366 = 4'he == w_addr_s1_0 | _GEN_3646; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6367 = 4'hf == w_addr_s1_0 | _GEN_3647; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6368 = wen_35 ? _GEN_6336 : data_0_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6369 = wen_35 ? _GEN_6337 : data_1_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6370 = wen_35 ? _GEN_6338 : data_2_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6371 = wen_35 ? _GEN_6339 : data_3_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6372 = wen_35 ? _GEN_6340 : data_4_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6373 = wen_35 ? _GEN_6341 : data_5_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6374 = wen_35 ? _GEN_6342 : data_6_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6375 = wen_35 ? _GEN_6343 : data_7_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6376 = wen_35 ? _GEN_6344 : data_8_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6377 = wen_35 ? _GEN_6345 : data_9_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6378 = wen_35 ? _GEN_6346 : data_10_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6379 = wen_35 ? _GEN_6347 : data_11_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6380 = wen_35 ? _GEN_6348 : data_12_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6381 = wen_35 ? _GEN_6349 : data_13_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6382 = wen_35 ? _GEN_6350 : data_14_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6383 = wen_35 ? _GEN_6351 : data_15_4_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6384 = wen_35 ? _GEN_6352 : _GEN_3632; // @[Sbuffer.scala 160:18]
  wire  _GEN_6385 = wen_35 ? _GEN_6353 : _GEN_3633; // @[Sbuffer.scala 160:18]
  wire  _GEN_6386 = wen_35 ? _GEN_6354 : _GEN_3634; // @[Sbuffer.scala 160:18]
  wire  _GEN_6387 = wen_35 ? _GEN_6355 : _GEN_3635; // @[Sbuffer.scala 160:18]
  wire  _GEN_6388 = wen_35 ? _GEN_6356 : _GEN_3636; // @[Sbuffer.scala 160:18]
  wire  _GEN_6389 = wen_35 ? _GEN_6357 : _GEN_3637; // @[Sbuffer.scala 160:18]
  wire  _GEN_6390 = wen_35 ? _GEN_6358 : _GEN_3638; // @[Sbuffer.scala 160:18]
  wire  _GEN_6391 = wen_35 ? _GEN_6359 : _GEN_3639; // @[Sbuffer.scala 160:18]
  wire  _GEN_6392 = wen_35 ? _GEN_6360 : _GEN_3640; // @[Sbuffer.scala 160:18]
  wire  _GEN_6393 = wen_35 ? _GEN_6361 : _GEN_3641; // @[Sbuffer.scala 160:18]
  wire  _GEN_6394 = wen_35 ? _GEN_6362 : _GEN_3642; // @[Sbuffer.scala 160:18]
  wire  _GEN_6395 = wen_35 ? _GEN_6363 : _GEN_3643; // @[Sbuffer.scala 160:18]
  wire  _GEN_6396 = wen_35 ? _GEN_6364 : _GEN_3644; // @[Sbuffer.scala 160:18]
  wire  _GEN_6397 = wen_35 ? _GEN_6365 : _GEN_3645; // @[Sbuffer.scala 160:18]
  wire  _GEN_6398 = wen_35 ? _GEN_6366 : _GEN_3646; // @[Sbuffer.scala 160:18]
  wire  _GEN_6399 = wen_35 ? _GEN_6367 : _GEN_3647; // @[Sbuffer.scala 160:18]
  wire  _wen_T_147 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_36 = w_valid_s1_0 & _wen_T_147; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6400 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6401 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6402 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6403 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6404 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6405 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6406 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6407 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6408 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6409 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6410 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6411 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6412 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6413 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6414 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6415 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_4_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6416 = 4'h0 == w_addr_s1_0 | _GEN_3648; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6417 = 4'h1 == w_addr_s1_0 | _GEN_3649; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6418 = 4'h2 == w_addr_s1_0 | _GEN_3650; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6419 = 4'h3 == w_addr_s1_0 | _GEN_3651; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6420 = 4'h4 == w_addr_s1_0 | _GEN_3652; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6421 = 4'h5 == w_addr_s1_0 | _GEN_3653; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6422 = 4'h6 == w_addr_s1_0 | _GEN_3654; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6423 = 4'h7 == w_addr_s1_0 | _GEN_3655; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6424 = 4'h8 == w_addr_s1_0 | _GEN_3656; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6425 = 4'h9 == w_addr_s1_0 | _GEN_3657; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6426 = 4'ha == w_addr_s1_0 | _GEN_3658; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6427 = 4'hb == w_addr_s1_0 | _GEN_3659; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6428 = 4'hc == w_addr_s1_0 | _GEN_3660; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6429 = 4'hd == w_addr_s1_0 | _GEN_3661; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6430 = 4'he == w_addr_s1_0 | _GEN_3662; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6431 = 4'hf == w_addr_s1_0 | _GEN_3663; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6432 = wen_36 ? _GEN_6400 : data_0_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6433 = wen_36 ? _GEN_6401 : data_1_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6434 = wen_36 ? _GEN_6402 : data_2_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6435 = wen_36 ? _GEN_6403 : data_3_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6436 = wen_36 ? _GEN_6404 : data_4_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6437 = wen_36 ? _GEN_6405 : data_5_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6438 = wen_36 ? _GEN_6406 : data_6_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6439 = wen_36 ? _GEN_6407 : data_7_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6440 = wen_36 ? _GEN_6408 : data_8_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6441 = wen_36 ? _GEN_6409 : data_9_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6442 = wen_36 ? _GEN_6410 : data_10_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6443 = wen_36 ? _GEN_6411 : data_11_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6444 = wen_36 ? _GEN_6412 : data_12_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6445 = wen_36 ? _GEN_6413 : data_13_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6446 = wen_36 ? _GEN_6414 : data_14_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6447 = wen_36 ? _GEN_6415 : data_15_4_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6448 = wen_36 ? _GEN_6416 : _GEN_3648; // @[Sbuffer.scala 160:18]
  wire  _GEN_6449 = wen_36 ? _GEN_6417 : _GEN_3649; // @[Sbuffer.scala 160:18]
  wire  _GEN_6450 = wen_36 ? _GEN_6418 : _GEN_3650; // @[Sbuffer.scala 160:18]
  wire  _GEN_6451 = wen_36 ? _GEN_6419 : _GEN_3651; // @[Sbuffer.scala 160:18]
  wire  _GEN_6452 = wen_36 ? _GEN_6420 : _GEN_3652; // @[Sbuffer.scala 160:18]
  wire  _GEN_6453 = wen_36 ? _GEN_6421 : _GEN_3653; // @[Sbuffer.scala 160:18]
  wire  _GEN_6454 = wen_36 ? _GEN_6422 : _GEN_3654; // @[Sbuffer.scala 160:18]
  wire  _GEN_6455 = wen_36 ? _GEN_6423 : _GEN_3655; // @[Sbuffer.scala 160:18]
  wire  _GEN_6456 = wen_36 ? _GEN_6424 : _GEN_3656; // @[Sbuffer.scala 160:18]
  wire  _GEN_6457 = wen_36 ? _GEN_6425 : _GEN_3657; // @[Sbuffer.scala 160:18]
  wire  _GEN_6458 = wen_36 ? _GEN_6426 : _GEN_3658; // @[Sbuffer.scala 160:18]
  wire  _GEN_6459 = wen_36 ? _GEN_6427 : _GEN_3659; // @[Sbuffer.scala 160:18]
  wire  _GEN_6460 = wen_36 ? _GEN_6428 : _GEN_3660; // @[Sbuffer.scala 160:18]
  wire  _GEN_6461 = wen_36 ? _GEN_6429 : _GEN_3661; // @[Sbuffer.scala 160:18]
  wire  _GEN_6462 = wen_36 ? _GEN_6430 : _GEN_3662; // @[Sbuffer.scala 160:18]
  wire  _GEN_6463 = wen_36 ? _GEN_6431 : _GEN_3663; // @[Sbuffer.scala 160:18]
  wire  _wen_T_151 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_37 = w_valid_s1_0 & _wen_T_151; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6464 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6465 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6466 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6467 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6468 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6469 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6470 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6471 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6472 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6473 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6474 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6475 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6476 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6477 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6478 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6479 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_4_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6480 = 4'h0 == w_addr_s1_0 | _GEN_3664; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6481 = 4'h1 == w_addr_s1_0 | _GEN_3665; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6482 = 4'h2 == w_addr_s1_0 | _GEN_3666; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6483 = 4'h3 == w_addr_s1_0 | _GEN_3667; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6484 = 4'h4 == w_addr_s1_0 | _GEN_3668; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6485 = 4'h5 == w_addr_s1_0 | _GEN_3669; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6486 = 4'h6 == w_addr_s1_0 | _GEN_3670; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6487 = 4'h7 == w_addr_s1_0 | _GEN_3671; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6488 = 4'h8 == w_addr_s1_0 | _GEN_3672; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6489 = 4'h9 == w_addr_s1_0 | _GEN_3673; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6490 = 4'ha == w_addr_s1_0 | _GEN_3674; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6491 = 4'hb == w_addr_s1_0 | _GEN_3675; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6492 = 4'hc == w_addr_s1_0 | _GEN_3676; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6493 = 4'hd == w_addr_s1_0 | _GEN_3677; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6494 = 4'he == w_addr_s1_0 | _GEN_3678; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6495 = 4'hf == w_addr_s1_0 | _GEN_3679; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6496 = wen_37 ? _GEN_6464 : data_0_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6497 = wen_37 ? _GEN_6465 : data_1_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6498 = wen_37 ? _GEN_6466 : data_2_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6499 = wen_37 ? _GEN_6467 : data_3_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6500 = wen_37 ? _GEN_6468 : data_4_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6501 = wen_37 ? _GEN_6469 : data_5_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6502 = wen_37 ? _GEN_6470 : data_6_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6503 = wen_37 ? _GEN_6471 : data_7_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6504 = wen_37 ? _GEN_6472 : data_8_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6505 = wen_37 ? _GEN_6473 : data_9_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6506 = wen_37 ? _GEN_6474 : data_10_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6507 = wen_37 ? _GEN_6475 : data_11_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6508 = wen_37 ? _GEN_6476 : data_12_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6509 = wen_37 ? _GEN_6477 : data_13_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6510 = wen_37 ? _GEN_6478 : data_14_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6511 = wen_37 ? _GEN_6479 : data_15_4_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6512 = wen_37 ? _GEN_6480 : _GEN_3664; // @[Sbuffer.scala 160:18]
  wire  _GEN_6513 = wen_37 ? _GEN_6481 : _GEN_3665; // @[Sbuffer.scala 160:18]
  wire  _GEN_6514 = wen_37 ? _GEN_6482 : _GEN_3666; // @[Sbuffer.scala 160:18]
  wire  _GEN_6515 = wen_37 ? _GEN_6483 : _GEN_3667; // @[Sbuffer.scala 160:18]
  wire  _GEN_6516 = wen_37 ? _GEN_6484 : _GEN_3668; // @[Sbuffer.scala 160:18]
  wire  _GEN_6517 = wen_37 ? _GEN_6485 : _GEN_3669; // @[Sbuffer.scala 160:18]
  wire  _GEN_6518 = wen_37 ? _GEN_6486 : _GEN_3670; // @[Sbuffer.scala 160:18]
  wire  _GEN_6519 = wen_37 ? _GEN_6487 : _GEN_3671; // @[Sbuffer.scala 160:18]
  wire  _GEN_6520 = wen_37 ? _GEN_6488 : _GEN_3672; // @[Sbuffer.scala 160:18]
  wire  _GEN_6521 = wen_37 ? _GEN_6489 : _GEN_3673; // @[Sbuffer.scala 160:18]
  wire  _GEN_6522 = wen_37 ? _GEN_6490 : _GEN_3674; // @[Sbuffer.scala 160:18]
  wire  _GEN_6523 = wen_37 ? _GEN_6491 : _GEN_3675; // @[Sbuffer.scala 160:18]
  wire  _GEN_6524 = wen_37 ? _GEN_6492 : _GEN_3676; // @[Sbuffer.scala 160:18]
  wire  _GEN_6525 = wen_37 ? _GEN_6493 : _GEN_3677; // @[Sbuffer.scala 160:18]
  wire  _GEN_6526 = wen_37 ? _GEN_6494 : _GEN_3678; // @[Sbuffer.scala 160:18]
  wire  _GEN_6527 = wen_37 ? _GEN_6495 : _GEN_3679; // @[Sbuffer.scala 160:18]
  wire  _wen_T_155 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_38 = w_valid_s1_0 & _wen_T_155; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6528 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6529 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6530 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6531 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6532 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6533 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6534 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6535 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6536 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6537 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6538 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6539 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6540 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6541 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6542 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6543 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_4_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6544 = 4'h0 == w_addr_s1_0 | _GEN_3680; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6545 = 4'h1 == w_addr_s1_0 | _GEN_3681; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6546 = 4'h2 == w_addr_s1_0 | _GEN_3682; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6547 = 4'h3 == w_addr_s1_0 | _GEN_3683; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6548 = 4'h4 == w_addr_s1_0 | _GEN_3684; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6549 = 4'h5 == w_addr_s1_0 | _GEN_3685; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6550 = 4'h6 == w_addr_s1_0 | _GEN_3686; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6551 = 4'h7 == w_addr_s1_0 | _GEN_3687; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6552 = 4'h8 == w_addr_s1_0 | _GEN_3688; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6553 = 4'h9 == w_addr_s1_0 | _GEN_3689; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6554 = 4'ha == w_addr_s1_0 | _GEN_3690; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6555 = 4'hb == w_addr_s1_0 | _GEN_3691; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6556 = 4'hc == w_addr_s1_0 | _GEN_3692; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6557 = 4'hd == w_addr_s1_0 | _GEN_3693; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6558 = 4'he == w_addr_s1_0 | _GEN_3694; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6559 = 4'hf == w_addr_s1_0 | _GEN_3695; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6560 = wen_38 ? _GEN_6528 : data_0_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6561 = wen_38 ? _GEN_6529 : data_1_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6562 = wen_38 ? _GEN_6530 : data_2_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6563 = wen_38 ? _GEN_6531 : data_3_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6564 = wen_38 ? _GEN_6532 : data_4_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6565 = wen_38 ? _GEN_6533 : data_5_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6566 = wen_38 ? _GEN_6534 : data_6_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6567 = wen_38 ? _GEN_6535 : data_7_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6568 = wen_38 ? _GEN_6536 : data_8_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6569 = wen_38 ? _GEN_6537 : data_9_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6570 = wen_38 ? _GEN_6538 : data_10_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6571 = wen_38 ? _GEN_6539 : data_11_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6572 = wen_38 ? _GEN_6540 : data_12_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6573 = wen_38 ? _GEN_6541 : data_13_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6574 = wen_38 ? _GEN_6542 : data_14_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6575 = wen_38 ? _GEN_6543 : data_15_4_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6576 = wen_38 ? _GEN_6544 : _GEN_3680; // @[Sbuffer.scala 160:18]
  wire  _GEN_6577 = wen_38 ? _GEN_6545 : _GEN_3681; // @[Sbuffer.scala 160:18]
  wire  _GEN_6578 = wen_38 ? _GEN_6546 : _GEN_3682; // @[Sbuffer.scala 160:18]
  wire  _GEN_6579 = wen_38 ? _GEN_6547 : _GEN_3683; // @[Sbuffer.scala 160:18]
  wire  _GEN_6580 = wen_38 ? _GEN_6548 : _GEN_3684; // @[Sbuffer.scala 160:18]
  wire  _GEN_6581 = wen_38 ? _GEN_6549 : _GEN_3685; // @[Sbuffer.scala 160:18]
  wire  _GEN_6582 = wen_38 ? _GEN_6550 : _GEN_3686; // @[Sbuffer.scala 160:18]
  wire  _GEN_6583 = wen_38 ? _GEN_6551 : _GEN_3687; // @[Sbuffer.scala 160:18]
  wire  _GEN_6584 = wen_38 ? _GEN_6552 : _GEN_3688; // @[Sbuffer.scala 160:18]
  wire  _GEN_6585 = wen_38 ? _GEN_6553 : _GEN_3689; // @[Sbuffer.scala 160:18]
  wire  _GEN_6586 = wen_38 ? _GEN_6554 : _GEN_3690; // @[Sbuffer.scala 160:18]
  wire  _GEN_6587 = wen_38 ? _GEN_6555 : _GEN_3691; // @[Sbuffer.scala 160:18]
  wire  _GEN_6588 = wen_38 ? _GEN_6556 : _GEN_3692; // @[Sbuffer.scala 160:18]
  wire  _GEN_6589 = wen_38 ? _GEN_6557 : _GEN_3693; // @[Sbuffer.scala 160:18]
  wire  _GEN_6590 = wen_38 ? _GEN_6558 : _GEN_3694; // @[Sbuffer.scala 160:18]
  wire  _GEN_6591 = wen_38 ? _GEN_6559 : _GEN_3695; // @[Sbuffer.scala 160:18]
  wire  _wen_T_159 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h4 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_39 = w_valid_s1_0 & _wen_T_159; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6592 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6593 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6594 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6595 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6596 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6597 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6598 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6599 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6600 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6601 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6602 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6603 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6604 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6605 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6606 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6607 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_4_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6608 = 4'h0 == w_addr_s1_0 | _GEN_3696; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6609 = 4'h1 == w_addr_s1_0 | _GEN_3697; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6610 = 4'h2 == w_addr_s1_0 | _GEN_3698; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6611 = 4'h3 == w_addr_s1_0 | _GEN_3699; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6612 = 4'h4 == w_addr_s1_0 | _GEN_3700; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6613 = 4'h5 == w_addr_s1_0 | _GEN_3701; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6614 = 4'h6 == w_addr_s1_0 | _GEN_3702; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6615 = 4'h7 == w_addr_s1_0 | _GEN_3703; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6616 = 4'h8 == w_addr_s1_0 | _GEN_3704; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6617 = 4'h9 == w_addr_s1_0 | _GEN_3705; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6618 = 4'ha == w_addr_s1_0 | _GEN_3706; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6619 = 4'hb == w_addr_s1_0 | _GEN_3707; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6620 = 4'hc == w_addr_s1_0 | _GEN_3708; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6621 = 4'hd == w_addr_s1_0 | _GEN_3709; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6622 = 4'he == w_addr_s1_0 | _GEN_3710; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6623 = 4'hf == w_addr_s1_0 | _GEN_3711; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6624 = wen_39 ? _GEN_6592 : data_0_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6625 = wen_39 ? _GEN_6593 : data_1_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6626 = wen_39 ? _GEN_6594 : data_2_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6627 = wen_39 ? _GEN_6595 : data_3_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6628 = wen_39 ? _GEN_6596 : data_4_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6629 = wen_39 ? _GEN_6597 : data_5_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6630 = wen_39 ? _GEN_6598 : data_6_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6631 = wen_39 ? _GEN_6599 : data_7_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6632 = wen_39 ? _GEN_6600 : data_8_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6633 = wen_39 ? _GEN_6601 : data_9_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6634 = wen_39 ? _GEN_6602 : data_10_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6635 = wen_39 ? _GEN_6603 : data_11_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6636 = wen_39 ? _GEN_6604 : data_12_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6637 = wen_39 ? _GEN_6605 : data_13_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6638 = wen_39 ? _GEN_6606 : data_14_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6639 = wen_39 ? _GEN_6607 : data_15_4_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6640 = wen_39 ? _GEN_6608 : _GEN_3696; // @[Sbuffer.scala 160:18]
  wire  _GEN_6641 = wen_39 ? _GEN_6609 : _GEN_3697; // @[Sbuffer.scala 160:18]
  wire  _GEN_6642 = wen_39 ? _GEN_6610 : _GEN_3698; // @[Sbuffer.scala 160:18]
  wire  _GEN_6643 = wen_39 ? _GEN_6611 : _GEN_3699; // @[Sbuffer.scala 160:18]
  wire  _GEN_6644 = wen_39 ? _GEN_6612 : _GEN_3700; // @[Sbuffer.scala 160:18]
  wire  _GEN_6645 = wen_39 ? _GEN_6613 : _GEN_3701; // @[Sbuffer.scala 160:18]
  wire  _GEN_6646 = wen_39 ? _GEN_6614 : _GEN_3702; // @[Sbuffer.scala 160:18]
  wire  _GEN_6647 = wen_39 ? _GEN_6615 : _GEN_3703; // @[Sbuffer.scala 160:18]
  wire  _GEN_6648 = wen_39 ? _GEN_6616 : _GEN_3704; // @[Sbuffer.scala 160:18]
  wire  _GEN_6649 = wen_39 ? _GEN_6617 : _GEN_3705; // @[Sbuffer.scala 160:18]
  wire  _GEN_6650 = wen_39 ? _GEN_6618 : _GEN_3706; // @[Sbuffer.scala 160:18]
  wire  _GEN_6651 = wen_39 ? _GEN_6619 : _GEN_3707; // @[Sbuffer.scala 160:18]
  wire  _GEN_6652 = wen_39 ? _GEN_6620 : _GEN_3708; // @[Sbuffer.scala 160:18]
  wire  _GEN_6653 = wen_39 ? _GEN_6621 : _GEN_3709; // @[Sbuffer.scala 160:18]
  wire  _GEN_6654 = wen_39 ? _GEN_6622 : _GEN_3710; // @[Sbuffer.scala 160:18]
  wire  _GEN_6655 = wen_39 ? _GEN_6623 : _GEN_3711; // @[Sbuffer.scala 160:18]
  wire  _wen_T_163 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_40 = w_valid_s1_0 & _wen_T_163; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6656 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6657 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6658 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6659 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6660 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6661 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6662 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6663 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6664 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6665 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6666 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6667 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6668 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6669 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6670 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6671 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_5_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6672 = 4'h0 == w_addr_s1_0 | _GEN_3712; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6673 = 4'h1 == w_addr_s1_0 | _GEN_3713; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6674 = 4'h2 == w_addr_s1_0 | _GEN_3714; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6675 = 4'h3 == w_addr_s1_0 | _GEN_3715; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6676 = 4'h4 == w_addr_s1_0 | _GEN_3716; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6677 = 4'h5 == w_addr_s1_0 | _GEN_3717; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6678 = 4'h6 == w_addr_s1_0 | _GEN_3718; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6679 = 4'h7 == w_addr_s1_0 | _GEN_3719; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6680 = 4'h8 == w_addr_s1_0 | _GEN_3720; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6681 = 4'h9 == w_addr_s1_0 | _GEN_3721; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6682 = 4'ha == w_addr_s1_0 | _GEN_3722; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6683 = 4'hb == w_addr_s1_0 | _GEN_3723; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6684 = 4'hc == w_addr_s1_0 | _GEN_3724; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6685 = 4'hd == w_addr_s1_0 | _GEN_3725; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6686 = 4'he == w_addr_s1_0 | _GEN_3726; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6687 = 4'hf == w_addr_s1_0 | _GEN_3727; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6688 = wen_40 ? _GEN_6656 : data_0_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6689 = wen_40 ? _GEN_6657 : data_1_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6690 = wen_40 ? _GEN_6658 : data_2_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6691 = wen_40 ? _GEN_6659 : data_3_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6692 = wen_40 ? _GEN_6660 : data_4_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6693 = wen_40 ? _GEN_6661 : data_5_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6694 = wen_40 ? _GEN_6662 : data_6_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6695 = wen_40 ? _GEN_6663 : data_7_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6696 = wen_40 ? _GEN_6664 : data_8_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6697 = wen_40 ? _GEN_6665 : data_9_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6698 = wen_40 ? _GEN_6666 : data_10_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6699 = wen_40 ? _GEN_6667 : data_11_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6700 = wen_40 ? _GEN_6668 : data_12_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6701 = wen_40 ? _GEN_6669 : data_13_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6702 = wen_40 ? _GEN_6670 : data_14_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6703 = wen_40 ? _GEN_6671 : data_15_5_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6704 = wen_40 ? _GEN_6672 : _GEN_3712; // @[Sbuffer.scala 160:18]
  wire  _GEN_6705 = wen_40 ? _GEN_6673 : _GEN_3713; // @[Sbuffer.scala 160:18]
  wire  _GEN_6706 = wen_40 ? _GEN_6674 : _GEN_3714; // @[Sbuffer.scala 160:18]
  wire  _GEN_6707 = wen_40 ? _GEN_6675 : _GEN_3715; // @[Sbuffer.scala 160:18]
  wire  _GEN_6708 = wen_40 ? _GEN_6676 : _GEN_3716; // @[Sbuffer.scala 160:18]
  wire  _GEN_6709 = wen_40 ? _GEN_6677 : _GEN_3717; // @[Sbuffer.scala 160:18]
  wire  _GEN_6710 = wen_40 ? _GEN_6678 : _GEN_3718; // @[Sbuffer.scala 160:18]
  wire  _GEN_6711 = wen_40 ? _GEN_6679 : _GEN_3719; // @[Sbuffer.scala 160:18]
  wire  _GEN_6712 = wen_40 ? _GEN_6680 : _GEN_3720; // @[Sbuffer.scala 160:18]
  wire  _GEN_6713 = wen_40 ? _GEN_6681 : _GEN_3721; // @[Sbuffer.scala 160:18]
  wire  _GEN_6714 = wen_40 ? _GEN_6682 : _GEN_3722; // @[Sbuffer.scala 160:18]
  wire  _GEN_6715 = wen_40 ? _GEN_6683 : _GEN_3723; // @[Sbuffer.scala 160:18]
  wire  _GEN_6716 = wen_40 ? _GEN_6684 : _GEN_3724; // @[Sbuffer.scala 160:18]
  wire  _GEN_6717 = wen_40 ? _GEN_6685 : _GEN_3725; // @[Sbuffer.scala 160:18]
  wire  _GEN_6718 = wen_40 ? _GEN_6686 : _GEN_3726; // @[Sbuffer.scala 160:18]
  wire  _GEN_6719 = wen_40 ? _GEN_6687 : _GEN_3727; // @[Sbuffer.scala 160:18]
  wire  _wen_T_167 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_41 = w_valid_s1_0 & _wen_T_167; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6720 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6721 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6722 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6723 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6724 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6725 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6726 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6727 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6728 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6729 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6730 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6731 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6732 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6733 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6734 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6735 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_5_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6736 = 4'h0 == w_addr_s1_0 | _GEN_3728; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6737 = 4'h1 == w_addr_s1_0 | _GEN_3729; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6738 = 4'h2 == w_addr_s1_0 | _GEN_3730; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6739 = 4'h3 == w_addr_s1_0 | _GEN_3731; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6740 = 4'h4 == w_addr_s1_0 | _GEN_3732; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6741 = 4'h5 == w_addr_s1_0 | _GEN_3733; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6742 = 4'h6 == w_addr_s1_0 | _GEN_3734; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6743 = 4'h7 == w_addr_s1_0 | _GEN_3735; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6744 = 4'h8 == w_addr_s1_0 | _GEN_3736; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6745 = 4'h9 == w_addr_s1_0 | _GEN_3737; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6746 = 4'ha == w_addr_s1_0 | _GEN_3738; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6747 = 4'hb == w_addr_s1_0 | _GEN_3739; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6748 = 4'hc == w_addr_s1_0 | _GEN_3740; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6749 = 4'hd == w_addr_s1_0 | _GEN_3741; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6750 = 4'he == w_addr_s1_0 | _GEN_3742; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6751 = 4'hf == w_addr_s1_0 | _GEN_3743; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6752 = wen_41 ? _GEN_6720 : data_0_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6753 = wen_41 ? _GEN_6721 : data_1_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6754 = wen_41 ? _GEN_6722 : data_2_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6755 = wen_41 ? _GEN_6723 : data_3_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6756 = wen_41 ? _GEN_6724 : data_4_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6757 = wen_41 ? _GEN_6725 : data_5_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6758 = wen_41 ? _GEN_6726 : data_6_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6759 = wen_41 ? _GEN_6727 : data_7_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6760 = wen_41 ? _GEN_6728 : data_8_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6761 = wen_41 ? _GEN_6729 : data_9_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6762 = wen_41 ? _GEN_6730 : data_10_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6763 = wen_41 ? _GEN_6731 : data_11_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6764 = wen_41 ? _GEN_6732 : data_12_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6765 = wen_41 ? _GEN_6733 : data_13_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6766 = wen_41 ? _GEN_6734 : data_14_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6767 = wen_41 ? _GEN_6735 : data_15_5_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6768 = wen_41 ? _GEN_6736 : _GEN_3728; // @[Sbuffer.scala 160:18]
  wire  _GEN_6769 = wen_41 ? _GEN_6737 : _GEN_3729; // @[Sbuffer.scala 160:18]
  wire  _GEN_6770 = wen_41 ? _GEN_6738 : _GEN_3730; // @[Sbuffer.scala 160:18]
  wire  _GEN_6771 = wen_41 ? _GEN_6739 : _GEN_3731; // @[Sbuffer.scala 160:18]
  wire  _GEN_6772 = wen_41 ? _GEN_6740 : _GEN_3732; // @[Sbuffer.scala 160:18]
  wire  _GEN_6773 = wen_41 ? _GEN_6741 : _GEN_3733; // @[Sbuffer.scala 160:18]
  wire  _GEN_6774 = wen_41 ? _GEN_6742 : _GEN_3734; // @[Sbuffer.scala 160:18]
  wire  _GEN_6775 = wen_41 ? _GEN_6743 : _GEN_3735; // @[Sbuffer.scala 160:18]
  wire  _GEN_6776 = wen_41 ? _GEN_6744 : _GEN_3736; // @[Sbuffer.scala 160:18]
  wire  _GEN_6777 = wen_41 ? _GEN_6745 : _GEN_3737; // @[Sbuffer.scala 160:18]
  wire  _GEN_6778 = wen_41 ? _GEN_6746 : _GEN_3738; // @[Sbuffer.scala 160:18]
  wire  _GEN_6779 = wen_41 ? _GEN_6747 : _GEN_3739; // @[Sbuffer.scala 160:18]
  wire  _GEN_6780 = wen_41 ? _GEN_6748 : _GEN_3740; // @[Sbuffer.scala 160:18]
  wire  _GEN_6781 = wen_41 ? _GEN_6749 : _GEN_3741; // @[Sbuffer.scala 160:18]
  wire  _GEN_6782 = wen_41 ? _GEN_6750 : _GEN_3742; // @[Sbuffer.scala 160:18]
  wire  _GEN_6783 = wen_41 ? _GEN_6751 : _GEN_3743; // @[Sbuffer.scala 160:18]
  wire  _wen_T_171 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_42 = w_valid_s1_0 & _wen_T_171; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6784 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6785 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6786 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6787 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6788 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6789 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6790 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6791 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6792 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6793 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6794 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6795 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6796 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6797 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6798 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6799 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_5_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6800 = 4'h0 == w_addr_s1_0 | _GEN_3744; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6801 = 4'h1 == w_addr_s1_0 | _GEN_3745; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6802 = 4'h2 == w_addr_s1_0 | _GEN_3746; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6803 = 4'h3 == w_addr_s1_0 | _GEN_3747; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6804 = 4'h4 == w_addr_s1_0 | _GEN_3748; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6805 = 4'h5 == w_addr_s1_0 | _GEN_3749; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6806 = 4'h6 == w_addr_s1_0 | _GEN_3750; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6807 = 4'h7 == w_addr_s1_0 | _GEN_3751; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6808 = 4'h8 == w_addr_s1_0 | _GEN_3752; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6809 = 4'h9 == w_addr_s1_0 | _GEN_3753; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6810 = 4'ha == w_addr_s1_0 | _GEN_3754; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6811 = 4'hb == w_addr_s1_0 | _GEN_3755; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6812 = 4'hc == w_addr_s1_0 | _GEN_3756; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6813 = 4'hd == w_addr_s1_0 | _GEN_3757; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6814 = 4'he == w_addr_s1_0 | _GEN_3758; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6815 = 4'hf == w_addr_s1_0 | _GEN_3759; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6816 = wen_42 ? _GEN_6784 : data_0_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6817 = wen_42 ? _GEN_6785 : data_1_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6818 = wen_42 ? _GEN_6786 : data_2_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6819 = wen_42 ? _GEN_6787 : data_3_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6820 = wen_42 ? _GEN_6788 : data_4_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6821 = wen_42 ? _GEN_6789 : data_5_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6822 = wen_42 ? _GEN_6790 : data_6_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6823 = wen_42 ? _GEN_6791 : data_7_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6824 = wen_42 ? _GEN_6792 : data_8_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6825 = wen_42 ? _GEN_6793 : data_9_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6826 = wen_42 ? _GEN_6794 : data_10_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6827 = wen_42 ? _GEN_6795 : data_11_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6828 = wen_42 ? _GEN_6796 : data_12_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6829 = wen_42 ? _GEN_6797 : data_13_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6830 = wen_42 ? _GEN_6798 : data_14_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6831 = wen_42 ? _GEN_6799 : data_15_5_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6832 = wen_42 ? _GEN_6800 : _GEN_3744; // @[Sbuffer.scala 160:18]
  wire  _GEN_6833 = wen_42 ? _GEN_6801 : _GEN_3745; // @[Sbuffer.scala 160:18]
  wire  _GEN_6834 = wen_42 ? _GEN_6802 : _GEN_3746; // @[Sbuffer.scala 160:18]
  wire  _GEN_6835 = wen_42 ? _GEN_6803 : _GEN_3747; // @[Sbuffer.scala 160:18]
  wire  _GEN_6836 = wen_42 ? _GEN_6804 : _GEN_3748; // @[Sbuffer.scala 160:18]
  wire  _GEN_6837 = wen_42 ? _GEN_6805 : _GEN_3749; // @[Sbuffer.scala 160:18]
  wire  _GEN_6838 = wen_42 ? _GEN_6806 : _GEN_3750; // @[Sbuffer.scala 160:18]
  wire  _GEN_6839 = wen_42 ? _GEN_6807 : _GEN_3751; // @[Sbuffer.scala 160:18]
  wire  _GEN_6840 = wen_42 ? _GEN_6808 : _GEN_3752; // @[Sbuffer.scala 160:18]
  wire  _GEN_6841 = wen_42 ? _GEN_6809 : _GEN_3753; // @[Sbuffer.scala 160:18]
  wire  _GEN_6842 = wen_42 ? _GEN_6810 : _GEN_3754; // @[Sbuffer.scala 160:18]
  wire  _GEN_6843 = wen_42 ? _GEN_6811 : _GEN_3755; // @[Sbuffer.scala 160:18]
  wire  _GEN_6844 = wen_42 ? _GEN_6812 : _GEN_3756; // @[Sbuffer.scala 160:18]
  wire  _GEN_6845 = wen_42 ? _GEN_6813 : _GEN_3757; // @[Sbuffer.scala 160:18]
  wire  _GEN_6846 = wen_42 ? _GEN_6814 : _GEN_3758; // @[Sbuffer.scala 160:18]
  wire  _GEN_6847 = wen_42 ? _GEN_6815 : _GEN_3759; // @[Sbuffer.scala 160:18]
  wire  _wen_T_175 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_43 = w_valid_s1_0 & _wen_T_175; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6848 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6849 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6850 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6851 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6852 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6853 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6854 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6855 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6856 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6857 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6858 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6859 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6860 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6861 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6862 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6863 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_5_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6864 = 4'h0 == w_addr_s1_0 | _GEN_3760; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6865 = 4'h1 == w_addr_s1_0 | _GEN_3761; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6866 = 4'h2 == w_addr_s1_0 | _GEN_3762; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6867 = 4'h3 == w_addr_s1_0 | _GEN_3763; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6868 = 4'h4 == w_addr_s1_0 | _GEN_3764; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6869 = 4'h5 == w_addr_s1_0 | _GEN_3765; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6870 = 4'h6 == w_addr_s1_0 | _GEN_3766; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6871 = 4'h7 == w_addr_s1_0 | _GEN_3767; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6872 = 4'h8 == w_addr_s1_0 | _GEN_3768; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6873 = 4'h9 == w_addr_s1_0 | _GEN_3769; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6874 = 4'ha == w_addr_s1_0 | _GEN_3770; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6875 = 4'hb == w_addr_s1_0 | _GEN_3771; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6876 = 4'hc == w_addr_s1_0 | _GEN_3772; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6877 = 4'hd == w_addr_s1_0 | _GEN_3773; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6878 = 4'he == w_addr_s1_0 | _GEN_3774; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6879 = 4'hf == w_addr_s1_0 | _GEN_3775; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6880 = wen_43 ? _GEN_6848 : data_0_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6881 = wen_43 ? _GEN_6849 : data_1_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6882 = wen_43 ? _GEN_6850 : data_2_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6883 = wen_43 ? _GEN_6851 : data_3_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6884 = wen_43 ? _GEN_6852 : data_4_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6885 = wen_43 ? _GEN_6853 : data_5_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6886 = wen_43 ? _GEN_6854 : data_6_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6887 = wen_43 ? _GEN_6855 : data_7_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6888 = wen_43 ? _GEN_6856 : data_8_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6889 = wen_43 ? _GEN_6857 : data_9_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6890 = wen_43 ? _GEN_6858 : data_10_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6891 = wen_43 ? _GEN_6859 : data_11_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6892 = wen_43 ? _GEN_6860 : data_12_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6893 = wen_43 ? _GEN_6861 : data_13_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6894 = wen_43 ? _GEN_6862 : data_14_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6895 = wen_43 ? _GEN_6863 : data_15_5_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6896 = wen_43 ? _GEN_6864 : _GEN_3760; // @[Sbuffer.scala 160:18]
  wire  _GEN_6897 = wen_43 ? _GEN_6865 : _GEN_3761; // @[Sbuffer.scala 160:18]
  wire  _GEN_6898 = wen_43 ? _GEN_6866 : _GEN_3762; // @[Sbuffer.scala 160:18]
  wire  _GEN_6899 = wen_43 ? _GEN_6867 : _GEN_3763; // @[Sbuffer.scala 160:18]
  wire  _GEN_6900 = wen_43 ? _GEN_6868 : _GEN_3764; // @[Sbuffer.scala 160:18]
  wire  _GEN_6901 = wen_43 ? _GEN_6869 : _GEN_3765; // @[Sbuffer.scala 160:18]
  wire  _GEN_6902 = wen_43 ? _GEN_6870 : _GEN_3766; // @[Sbuffer.scala 160:18]
  wire  _GEN_6903 = wen_43 ? _GEN_6871 : _GEN_3767; // @[Sbuffer.scala 160:18]
  wire  _GEN_6904 = wen_43 ? _GEN_6872 : _GEN_3768; // @[Sbuffer.scala 160:18]
  wire  _GEN_6905 = wen_43 ? _GEN_6873 : _GEN_3769; // @[Sbuffer.scala 160:18]
  wire  _GEN_6906 = wen_43 ? _GEN_6874 : _GEN_3770; // @[Sbuffer.scala 160:18]
  wire  _GEN_6907 = wen_43 ? _GEN_6875 : _GEN_3771; // @[Sbuffer.scala 160:18]
  wire  _GEN_6908 = wen_43 ? _GEN_6876 : _GEN_3772; // @[Sbuffer.scala 160:18]
  wire  _GEN_6909 = wen_43 ? _GEN_6877 : _GEN_3773; // @[Sbuffer.scala 160:18]
  wire  _GEN_6910 = wen_43 ? _GEN_6878 : _GEN_3774; // @[Sbuffer.scala 160:18]
  wire  _GEN_6911 = wen_43 ? _GEN_6879 : _GEN_3775; // @[Sbuffer.scala 160:18]
  wire  _wen_T_179 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_44 = w_valid_s1_0 & _wen_T_179; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6912 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6913 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6914 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6915 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6916 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6917 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6918 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6919 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6920 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6921 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6922 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6923 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6924 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6925 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6926 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6927 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_5_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6928 = 4'h0 == w_addr_s1_0 | _GEN_3776; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6929 = 4'h1 == w_addr_s1_0 | _GEN_3777; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6930 = 4'h2 == w_addr_s1_0 | _GEN_3778; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6931 = 4'h3 == w_addr_s1_0 | _GEN_3779; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6932 = 4'h4 == w_addr_s1_0 | _GEN_3780; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6933 = 4'h5 == w_addr_s1_0 | _GEN_3781; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6934 = 4'h6 == w_addr_s1_0 | _GEN_3782; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6935 = 4'h7 == w_addr_s1_0 | _GEN_3783; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6936 = 4'h8 == w_addr_s1_0 | _GEN_3784; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6937 = 4'h9 == w_addr_s1_0 | _GEN_3785; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6938 = 4'ha == w_addr_s1_0 | _GEN_3786; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6939 = 4'hb == w_addr_s1_0 | _GEN_3787; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6940 = 4'hc == w_addr_s1_0 | _GEN_3788; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6941 = 4'hd == w_addr_s1_0 | _GEN_3789; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6942 = 4'he == w_addr_s1_0 | _GEN_3790; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6943 = 4'hf == w_addr_s1_0 | _GEN_3791; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_6944 = wen_44 ? _GEN_6912 : data_0_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6945 = wen_44 ? _GEN_6913 : data_1_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6946 = wen_44 ? _GEN_6914 : data_2_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6947 = wen_44 ? _GEN_6915 : data_3_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6948 = wen_44 ? _GEN_6916 : data_4_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6949 = wen_44 ? _GEN_6917 : data_5_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6950 = wen_44 ? _GEN_6918 : data_6_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6951 = wen_44 ? _GEN_6919 : data_7_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6952 = wen_44 ? _GEN_6920 : data_8_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6953 = wen_44 ? _GEN_6921 : data_9_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6954 = wen_44 ? _GEN_6922 : data_10_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6955 = wen_44 ? _GEN_6923 : data_11_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6956 = wen_44 ? _GEN_6924 : data_12_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6957 = wen_44 ? _GEN_6925 : data_13_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6958 = wen_44 ? _GEN_6926 : data_14_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_6959 = wen_44 ? _GEN_6927 : data_15_5_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_6960 = wen_44 ? _GEN_6928 : _GEN_3776; // @[Sbuffer.scala 160:18]
  wire  _GEN_6961 = wen_44 ? _GEN_6929 : _GEN_3777; // @[Sbuffer.scala 160:18]
  wire  _GEN_6962 = wen_44 ? _GEN_6930 : _GEN_3778; // @[Sbuffer.scala 160:18]
  wire  _GEN_6963 = wen_44 ? _GEN_6931 : _GEN_3779; // @[Sbuffer.scala 160:18]
  wire  _GEN_6964 = wen_44 ? _GEN_6932 : _GEN_3780; // @[Sbuffer.scala 160:18]
  wire  _GEN_6965 = wen_44 ? _GEN_6933 : _GEN_3781; // @[Sbuffer.scala 160:18]
  wire  _GEN_6966 = wen_44 ? _GEN_6934 : _GEN_3782; // @[Sbuffer.scala 160:18]
  wire  _GEN_6967 = wen_44 ? _GEN_6935 : _GEN_3783; // @[Sbuffer.scala 160:18]
  wire  _GEN_6968 = wen_44 ? _GEN_6936 : _GEN_3784; // @[Sbuffer.scala 160:18]
  wire  _GEN_6969 = wen_44 ? _GEN_6937 : _GEN_3785; // @[Sbuffer.scala 160:18]
  wire  _GEN_6970 = wen_44 ? _GEN_6938 : _GEN_3786; // @[Sbuffer.scala 160:18]
  wire  _GEN_6971 = wen_44 ? _GEN_6939 : _GEN_3787; // @[Sbuffer.scala 160:18]
  wire  _GEN_6972 = wen_44 ? _GEN_6940 : _GEN_3788; // @[Sbuffer.scala 160:18]
  wire  _GEN_6973 = wen_44 ? _GEN_6941 : _GEN_3789; // @[Sbuffer.scala 160:18]
  wire  _GEN_6974 = wen_44 ? _GEN_6942 : _GEN_3790; // @[Sbuffer.scala 160:18]
  wire  _GEN_6975 = wen_44 ? _GEN_6943 : _GEN_3791; // @[Sbuffer.scala 160:18]
  wire  _wen_T_183 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_45 = w_valid_s1_0 & _wen_T_183; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_6976 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6977 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6978 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6979 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6980 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6981 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6982 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6983 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6984 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6985 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6986 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6987 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6988 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6989 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6990 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_6991 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_5_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_6992 = 4'h0 == w_addr_s1_0 | _GEN_3792; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6993 = 4'h1 == w_addr_s1_0 | _GEN_3793; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6994 = 4'h2 == w_addr_s1_0 | _GEN_3794; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6995 = 4'h3 == w_addr_s1_0 | _GEN_3795; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6996 = 4'h4 == w_addr_s1_0 | _GEN_3796; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6997 = 4'h5 == w_addr_s1_0 | _GEN_3797; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6998 = 4'h6 == w_addr_s1_0 | _GEN_3798; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_6999 = 4'h7 == w_addr_s1_0 | _GEN_3799; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7000 = 4'h8 == w_addr_s1_0 | _GEN_3800; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7001 = 4'h9 == w_addr_s1_0 | _GEN_3801; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7002 = 4'ha == w_addr_s1_0 | _GEN_3802; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7003 = 4'hb == w_addr_s1_0 | _GEN_3803; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7004 = 4'hc == w_addr_s1_0 | _GEN_3804; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7005 = 4'hd == w_addr_s1_0 | _GEN_3805; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7006 = 4'he == w_addr_s1_0 | _GEN_3806; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7007 = 4'hf == w_addr_s1_0 | _GEN_3807; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7008 = wen_45 ? _GEN_6976 : data_0_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7009 = wen_45 ? _GEN_6977 : data_1_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7010 = wen_45 ? _GEN_6978 : data_2_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7011 = wen_45 ? _GEN_6979 : data_3_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7012 = wen_45 ? _GEN_6980 : data_4_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7013 = wen_45 ? _GEN_6981 : data_5_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7014 = wen_45 ? _GEN_6982 : data_6_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7015 = wen_45 ? _GEN_6983 : data_7_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7016 = wen_45 ? _GEN_6984 : data_8_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7017 = wen_45 ? _GEN_6985 : data_9_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7018 = wen_45 ? _GEN_6986 : data_10_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7019 = wen_45 ? _GEN_6987 : data_11_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7020 = wen_45 ? _GEN_6988 : data_12_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7021 = wen_45 ? _GEN_6989 : data_13_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7022 = wen_45 ? _GEN_6990 : data_14_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7023 = wen_45 ? _GEN_6991 : data_15_5_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7024 = wen_45 ? _GEN_6992 : _GEN_3792; // @[Sbuffer.scala 160:18]
  wire  _GEN_7025 = wen_45 ? _GEN_6993 : _GEN_3793; // @[Sbuffer.scala 160:18]
  wire  _GEN_7026 = wen_45 ? _GEN_6994 : _GEN_3794; // @[Sbuffer.scala 160:18]
  wire  _GEN_7027 = wen_45 ? _GEN_6995 : _GEN_3795; // @[Sbuffer.scala 160:18]
  wire  _GEN_7028 = wen_45 ? _GEN_6996 : _GEN_3796; // @[Sbuffer.scala 160:18]
  wire  _GEN_7029 = wen_45 ? _GEN_6997 : _GEN_3797; // @[Sbuffer.scala 160:18]
  wire  _GEN_7030 = wen_45 ? _GEN_6998 : _GEN_3798; // @[Sbuffer.scala 160:18]
  wire  _GEN_7031 = wen_45 ? _GEN_6999 : _GEN_3799; // @[Sbuffer.scala 160:18]
  wire  _GEN_7032 = wen_45 ? _GEN_7000 : _GEN_3800; // @[Sbuffer.scala 160:18]
  wire  _GEN_7033 = wen_45 ? _GEN_7001 : _GEN_3801; // @[Sbuffer.scala 160:18]
  wire  _GEN_7034 = wen_45 ? _GEN_7002 : _GEN_3802; // @[Sbuffer.scala 160:18]
  wire  _GEN_7035 = wen_45 ? _GEN_7003 : _GEN_3803; // @[Sbuffer.scala 160:18]
  wire  _GEN_7036 = wen_45 ? _GEN_7004 : _GEN_3804; // @[Sbuffer.scala 160:18]
  wire  _GEN_7037 = wen_45 ? _GEN_7005 : _GEN_3805; // @[Sbuffer.scala 160:18]
  wire  _GEN_7038 = wen_45 ? _GEN_7006 : _GEN_3806; // @[Sbuffer.scala 160:18]
  wire  _GEN_7039 = wen_45 ? _GEN_7007 : _GEN_3807; // @[Sbuffer.scala 160:18]
  wire  _wen_T_187 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_46 = w_valid_s1_0 & _wen_T_187; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7040 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7041 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7042 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7043 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7044 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7045 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7046 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7047 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7048 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7049 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7050 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7051 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7052 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7053 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7054 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7055 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_5_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7056 = 4'h0 == w_addr_s1_0 | _GEN_3808; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7057 = 4'h1 == w_addr_s1_0 | _GEN_3809; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7058 = 4'h2 == w_addr_s1_0 | _GEN_3810; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7059 = 4'h3 == w_addr_s1_0 | _GEN_3811; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7060 = 4'h4 == w_addr_s1_0 | _GEN_3812; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7061 = 4'h5 == w_addr_s1_0 | _GEN_3813; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7062 = 4'h6 == w_addr_s1_0 | _GEN_3814; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7063 = 4'h7 == w_addr_s1_0 | _GEN_3815; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7064 = 4'h8 == w_addr_s1_0 | _GEN_3816; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7065 = 4'h9 == w_addr_s1_0 | _GEN_3817; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7066 = 4'ha == w_addr_s1_0 | _GEN_3818; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7067 = 4'hb == w_addr_s1_0 | _GEN_3819; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7068 = 4'hc == w_addr_s1_0 | _GEN_3820; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7069 = 4'hd == w_addr_s1_0 | _GEN_3821; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7070 = 4'he == w_addr_s1_0 | _GEN_3822; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7071 = 4'hf == w_addr_s1_0 | _GEN_3823; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7072 = wen_46 ? _GEN_7040 : data_0_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7073 = wen_46 ? _GEN_7041 : data_1_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7074 = wen_46 ? _GEN_7042 : data_2_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7075 = wen_46 ? _GEN_7043 : data_3_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7076 = wen_46 ? _GEN_7044 : data_4_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7077 = wen_46 ? _GEN_7045 : data_5_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7078 = wen_46 ? _GEN_7046 : data_6_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7079 = wen_46 ? _GEN_7047 : data_7_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7080 = wen_46 ? _GEN_7048 : data_8_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7081 = wen_46 ? _GEN_7049 : data_9_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7082 = wen_46 ? _GEN_7050 : data_10_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7083 = wen_46 ? _GEN_7051 : data_11_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7084 = wen_46 ? _GEN_7052 : data_12_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7085 = wen_46 ? _GEN_7053 : data_13_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7086 = wen_46 ? _GEN_7054 : data_14_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7087 = wen_46 ? _GEN_7055 : data_15_5_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7088 = wen_46 ? _GEN_7056 : _GEN_3808; // @[Sbuffer.scala 160:18]
  wire  _GEN_7089 = wen_46 ? _GEN_7057 : _GEN_3809; // @[Sbuffer.scala 160:18]
  wire  _GEN_7090 = wen_46 ? _GEN_7058 : _GEN_3810; // @[Sbuffer.scala 160:18]
  wire  _GEN_7091 = wen_46 ? _GEN_7059 : _GEN_3811; // @[Sbuffer.scala 160:18]
  wire  _GEN_7092 = wen_46 ? _GEN_7060 : _GEN_3812; // @[Sbuffer.scala 160:18]
  wire  _GEN_7093 = wen_46 ? _GEN_7061 : _GEN_3813; // @[Sbuffer.scala 160:18]
  wire  _GEN_7094 = wen_46 ? _GEN_7062 : _GEN_3814; // @[Sbuffer.scala 160:18]
  wire  _GEN_7095 = wen_46 ? _GEN_7063 : _GEN_3815; // @[Sbuffer.scala 160:18]
  wire  _GEN_7096 = wen_46 ? _GEN_7064 : _GEN_3816; // @[Sbuffer.scala 160:18]
  wire  _GEN_7097 = wen_46 ? _GEN_7065 : _GEN_3817; // @[Sbuffer.scala 160:18]
  wire  _GEN_7098 = wen_46 ? _GEN_7066 : _GEN_3818; // @[Sbuffer.scala 160:18]
  wire  _GEN_7099 = wen_46 ? _GEN_7067 : _GEN_3819; // @[Sbuffer.scala 160:18]
  wire  _GEN_7100 = wen_46 ? _GEN_7068 : _GEN_3820; // @[Sbuffer.scala 160:18]
  wire  _GEN_7101 = wen_46 ? _GEN_7069 : _GEN_3821; // @[Sbuffer.scala 160:18]
  wire  _GEN_7102 = wen_46 ? _GEN_7070 : _GEN_3822; // @[Sbuffer.scala 160:18]
  wire  _GEN_7103 = wen_46 ? _GEN_7071 : _GEN_3823; // @[Sbuffer.scala 160:18]
  wire  _wen_T_191 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h5 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_47 = w_valid_s1_0 & _wen_T_191; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7104 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7105 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7106 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7107 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7108 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7109 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7110 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7111 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7112 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7113 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7114 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7115 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7116 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7117 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7118 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7119 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_5_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7120 = 4'h0 == w_addr_s1_0 | _GEN_3824; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7121 = 4'h1 == w_addr_s1_0 | _GEN_3825; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7122 = 4'h2 == w_addr_s1_0 | _GEN_3826; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7123 = 4'h3 == w_addr_s1_0 | _GEN_3827; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7124 = 4'h4 == w_addr_s1_0 | _GEN_3828; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7125 = 4'h5 == w_addr_s1_0 | _GEN_3829; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7126 = 4'h6 == w_addr_s1_0 | _GEN_3830; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7127 = 4'h7 == w_addr_s1_0 | _GEN_3831; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7128 = 4'h8 == w_addr_s1_0 | _GEN_3832; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7129 = 4'h9 == w_addr_s1_0 | _GEN_3833; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7130 = 4'ha == w_addr_s1_0 | _GEN_3834; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7131 = 4'hb == w_addr_s1_0 | _GEN_3835; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7132 = 4'hc == w_addr_s1_0 | _GEN_3836; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7133 = 4'hd == w_addr_s1_0 | _GEN_3837; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7134 = 4'he == w_addr_s1_0 | _GEN_3838; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7135 = 4'hf == w_addr_s1_0 | _GEN_3839; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7136 = wen_47 ? _GEN_7104 : data_0_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7137 = wen_47 ? _GEN_7105 : data_1_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7138 = wen_47 ? _GEN_7106 : data_2_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7139 = wen_47 ? _GEN_7107 : data_3_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7140 = wen_47 ? _GEN_7108 : data_4_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7141 = wen_47 ? _GEN_7109 : data_5_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7142 = wen_47 ? _GEN_7110 : data_6_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7143 = wen_47 ? _GEN_7111 : data_7_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7144 = wen_47 ? _GEN_7112 : data_8_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7145 = wen_47 ? _GEN_7113 : data_9_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7146 = wen_47 ? _GEN_7114 : data_10_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7147 = wen_47 ? _GEN_7115 : data_11_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7148 = wen_47 ? _GEN_7116 : data_12_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7149 = wen_47 ? _GEN_7117 : data_13_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7150 = wen_47 ? _GEN_7118 : data_14_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7151 = wen_47 ? _GEN_7119 : data_15_5_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7152 = wen_47 ? _GEN_7120 : _GEN_3824; // @[Sbuffer.scala 160:18]
  wire  _GEN_7153 = wen_47 ? _GEN_7121 : _GEN_3825; // @[Sbuffer.scala 160:18]
  wire  _GEN_7154 = wen_47 ? _GEN_7122 : _GEN_3826; // @[Sbuffer.scala 160:18]
  wire  _GEN_7155 = wen_47 ? _GEN_7123 : _GEN_3827; // @[Sbuffer.scala 160:18]
  wire  _GEN_7156 = wen_47 ? _GEN_7124 : _GEN_3828; // @[Sbuffer.scala 160:18]
  wire  _GEN_7157 = wen_47 ? _GEN_7125 : _GEN_3829; // @[Sbuffer.scala 160:18]
  wire  _GEN_7158 = wen_47 ? _GEN_7126 : _GEN_3830; // @[Sbuffer.scala 160:18]
  wire  _GEN_7159 = wen_47 ? _GEN_7127 : _GEN_3831; // @[Sbuffer.scala 160:18]
  wire  _GEN_7160 = wen_47 ? _GEN_7128 : _GEN_3832; // @[Sbuffer.scala 160:18]
  wire  _GEN_7161 = wen_47 ? _GEN_7129 : _GEN_3833; // @[Sbuffer.scala 160:18]
  wire  _GEN_7162 = wen_47 ? _GEN_7130 : _GEN_3834; // @[Sbuffer.scala 160:18]
  wire  _GEN_7163 = wen_47 ? _GEN_7131 : _GEN_3835; // @[Sbuffer.scala 160:18]
  wire  _GEN_7164 = wen_47 ? _GEN_7132 : _GEN_3836; // @[Sbuffer.scala 160:18]
  wire  _GEN_7165 = wen_47 ? _GEN_7133 : _GEN_3837; // @[Sbuffer.scala 160:18]
  wire  _GEN_7166 = wen_47 ? _GEN_7134 : _GEN_3838; // @[Sbuffer.scala 160:18]
  wire  _GEN_7167 = wen_47 ? _GEN_7135 : _GEN_3839; // @[Sbuffer.scala 160:18]
  wire  _wen_T_195 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_48 = w_valid_s1_0 & _wen_T_195; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7168 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7169 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7170 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7171 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7172 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7173 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7174 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7175 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7176 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7177 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7178 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7179 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7180 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7181 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7182 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7183 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_6_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7184 = 4'h0 == w_addr_s1_0 | _GEN_3840; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7185 = 4'h1 == w_addr_s1_0 | _GEN_3841; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7186 = 4'h2 == w_addr_s1_0 | _GEN_3842; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7187 = 4'h3 == w_addr_s1_0 | _GEN_3843; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7188 = 4'h4 == w_addr_s1_0 | _GEN_3844; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7189 = 4'h5 == w_addr_s1_0 | _GEN_3845; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7190 = 4'h6 == w_addr_s1_0 | _GEN_3846; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7191 = 4'h7 == w_addr_s1_0 | _GEN_3847; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7192 = 4'h8 == w_addr_s1_0 | _GEN_3848; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7193 = 4'h9 == w_addr_s1_0 | _GEN_3849; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7194 = 4'ha == w_addr_s1_0 | _GEN_3850; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7195 = 4'hb == w_addr_s1_0 | _GEN_3851; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7196 = 4'hc == w_addr_s1_0 | _GEN_3852; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7197 = 4'hd == w_addr_s1_0 | _GEN_3853; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7198 = 4'he == w_addr_s1_0 | _GEN_3854; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7199 = 4'hf == w_addr_s1_0 | _GEN_3855; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7200 = wen_48 ? _GEN_7168 : data_0_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7201 = wen_48 ? _GEN_7169 : data_1_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7202 = wen_48 ? _GEN_7170 : data_2_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7203 = wen_48 ? _GEN_7171 : data_3_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7204 = wen_48 ? _GEN_7172 : data_4_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7205 = wen_48 ? _GEN_7173 : data_5_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7206 = wen_48 ? _GEN_7174 : data_6_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7207 = wen_48 ? _GEN_7175 : data_7_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7208 = wen_48 ? _GEN_7176 : data_8_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7209 = wen_48 ? _GEN_7177 : data_9_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7210 = wen_48 ? _GEN_7178 : data_10_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7211 = wen_48 ? _GEN_7179 : data_11_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7212 = wen_48 ? _GEN_7180 : data_12_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7213 = wen_48 ? _GEN_7181 : data_13_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7214 = wen_48 ? _GEN_7182 : data_14_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7215 = wen_48 ? _GEN_7183 : data_15_6_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7216 = wen_48 ? _GEN_7184 : _GEN_3840; // @[Sbuffer.scala 160:18]
  wire  _GEN_7217 = wen_48 ? _GEN_7185 : _GEN_3841; // @[Sbuffer.scala 160:18]
  wire  _GEN_7218 = wen_48 ? _GEN_7186 : _GEN_3842; // @[Sbuffer.scala 160:18]
  wire  _GEN_7219 = wen_48 ? _GEN_7187 : _GEN_3843; // @[Sbuffer.scala 160:18]
  wire  _GEN_7220 = wen_48 ? _GEN_7188 : _GEN_3844; // @[Sbuffer.scala 160:18]
  wire  _GEN_7221 = wen_48 ? _GEN_7189 : _GEN_3845; // @[Sbuffer.scala 160:18]
  wire  _GEN_7222 = wen_48 ? _GEN_7190 : _GEN_3846; // @[Sbuffer.scala 160:18]
  wire  _GEN_7223 = wen_48 ? _GEN_7191 : _GEN_3847; // @[Sbuffer.scala 160:18]
  wire  _GEN_7224 = wen_48 ? _GEN_7192 : _GEN_3848; // @[Sbuffer.scala 160:18]
  wire  _GEN_7225 = wen_48 ? _GEN_7193 : _GEN_3849; // @[Sbuffer.scala 160:18]
  wire  _GEN_7226 = wen_48 ? _GEN_7194 : _GEN_3850; // @[Sbuffer.scala 160:18]
  wire  _GEN_7227 = wen_48 ? _GEN_7195 : _GEN_3851; // @[Sbuffer.scala 160:18]
  wire  _GEN_7228 = wen_48 ? _GEN_7196 : _GEN_3852; // @[Sbuffer.scala 160:18]
  wire  _GEN_7229 = wen_48 ? _GEN_7197 : _GEN_3853; // @[Sbuffer.scala 160:18]
  wire  _GEN_7230 = wen_48 ? _GEN_7198 : _GEN_3854; // @[Sbuffer.scala 160:18]
  wire  _GEN_7231 = wen_48 ? _GEN_7199 : _GEN_3855; // @[Sbuffer.scala 160:18]
  wire  _wen_T_199 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_49 = w_valid_s1_0 & _wen_T_199; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7232 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7233 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7234 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7235 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7236 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7237 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7238 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7239 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7240 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7241 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7242 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7243 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7244 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7245 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7246 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7247 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_6_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7248 = 4'h0 == w_addr_s1_0 | _GEN_3856; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7249 = 4'h1 == w_addr_s1_0 | _GEN_3857; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7250 = 4'h2 == w_addr_s1_0 | _GEN_3858; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7251 = 4'h3 == w_addr_s1_0 | _GEN_3859; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7252 = 4'h4 == w_addr_s1_0 | _GEN_3860; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7253 = 4'h5 == w_addr_s1_0 | _GEN_3861; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7254 = 4'h6 == w_addr_s1_0 | _GEN_3862; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7255 = 4'h7 == w_addr_s1_0 | _GEN_3863; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7256 = 4'h8 == w_addr_s1_0 | _GEN_3864; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7257 = 4'h9 == w_addr_s1_0 | _GEN_3865; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7258 = 4'ha == w_addr_s1_0 | _GEN_3866; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7259 = 4'hb == w_addr_s1_0 | _GEN_3867; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7260 = 4'hc == w_addr_s1_0 | _GEN_3868; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7261 = 4'hd == w_addr_s1_0 | _GEN_3869; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7262 = 4'he == w_addr_s1_0 | _GEN_3870; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7263 = 4'hf == w_addr_s1_0 | _GEN_3871; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7264 = wen_49 ? _GEN_7232 : data_0_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7265 = wen_49 ? _GEN_7233 : data_1_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7266 = wen_49 ? _GEN_7234 : data_2_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7267 = wen_49 ? _GEN_7235 : data_3_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7268 = wen_49 ? _GEN_7236 : data_4_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7269 = wen_49 ? _GEN_7237 : data_5_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7270 = wen_49 ? _GEN_7238 : data_6_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7271 = wen_49 ? _GEN_7239 : data_7_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7272 = wen_49 ? _GEN_7240 : data_8_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7273 = wen_49 ? _GEN_7241 : data_9_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7274 = wen_49 ? _GEN_7242 : data_10_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7275 = wen_49 ? _GEN_7243 : data_11_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7276 = wen_49 ? _GEN_7244 : data_12_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7277 = wen_49 ? _GEN_7245 : data_13_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7278 = wen_49 ? _GEN_7246 : data_14_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7279 = wen_49 ? _GEN_7247 : data_15_6_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7280 = wen_49 ? _GEN_7248 : _GEN_3856; // @[Sbuffer.scala 160:18]
  wire  _GEN_7281 = wen_49 ? _GEN_7249 : _GEN_3857; // @[Sbuffer.scala 160:18]
  wire  _GEN_7282 = wen_49 ? _GEN_7250 : _GEN_3858; // @[Sbuffer.scala 160:18]
  wire  _GEN_7283 = wen_49 ? _GEN_7251 : _GEN_3859; // @[Sbuffer.scala 160:18]
  wire  _GEN_7284 = wen_49 ? _GEN_7252 : _GEN_3860; // @[Sbuffer.scala 160:18]
  wire  _GEN_7285 = wen_49 ? _GEN_7253 : _GEN_3861; // @[Sbuffer.scala 160:18]
  wire  _GEN_7286 = wen_49 ? _GEN_7254 : _GEN_3862; // @[Sbuffer.scala 160:18]
  wire  _GEN_7287 = wen_49 ? _GEN_7255 : _GEN_3863; // @[Sbuffer.scala 160:18]
  wire  _GEN_7288 = wen_49 ? _GEN_7256 : _GEN_3864; // @[Sbuffer.scala 160:18]
  wire  _GEN_7289 = wen_49 ? _GEN_7257 : _GEN_3865; // @[Sbuffer.scala 160:18]
  wire  _GEN_7290 = wen_49 ? _GEN_7258 : _GEN_3866; // @[Sbuffer.scala 160:18]
  wire  _GEN_7291 = wen_49 ? _GEN_7259 : _GEN_3867; // @[Sbuffer.scala 160:18]
  wire  _GEN_7292 = wen_49 ? _GEN_7260 : _GEN_3868; // @[Sbuffer.scala 160:18]
  wire  _GEN_7293 = wen_49 ? _GEN_7261 : _GEN_3869; // @[Sbuffer.scala 160:18]
  wire  _GEN_7294 = wen_49 ? _GEN_7262 : _GEN_3870; // @[Sbuffer.scala 160:18]
  wire  _GEN_7295 = wen_49 ? _GEN_7263 : _GEN_3871; // @[Sbuffer.scala 160:18]
  wire  _wen_T_203 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_50 = w_valid_s1_0 & _wen_T_203; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7296 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7297 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7298 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7299 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7300 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7301 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7302 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7303 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7304 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7305 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7306 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7307 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7308 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7309 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7310 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7311 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_6_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7312 = 4'h0 == w_addr_s1_0 | _GEN_3872; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7313 = 4'h1 == w_addr_s1_0 | _GEN_3873; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7314 = 4'h2 == w_addr_s1_0 | _GEN_3874; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7315 = 4'h3 == w_addr_s1_0 | _GEN_3875; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7316 = 4'h4 == w_addr_s1_0 | _GEN_3876; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7317 = 4'h5 == w_addr_s1_0 | _GEN_3877; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7318 = 4'h6 == w_addr_s1_0 | _GEN_3878; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7319 = 4'h7 == w_addr_s1_0 | _GEN_3879; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7320 = 4'h8 == w_addr_s1_0 | _GEN_3880; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7321 = 4'h9 == w_addr_s1_0 | _GEN_3881; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7322 = 4'ha == w_addr_s1_0 | _GEN_3882; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7323 = 4'hb == w_addr_s1_0 | _GEN_3883; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7324 = 4'hc == w_addr_s1_0 | _GEN_3884; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7325 = 4'hd == w_addr_s1_0 | _GEN_3885; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7326 = 4'he == w_addr_s1_0 | _GEN_3886; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7327 = 4'hf == w_addr_s1_0 | _GEN_3887; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7328 = wen_50 ? _GEN_7296 : data_0_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7329 = wen_50 ? _GEN_7297 : data_1_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7330 = wen_50 ? _GEN_7298 : data_2_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7331 = wen_50 ? _GEN_7299 : data_3_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7332 = wen_50 ? _GEN_7300 : data_4_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7333 = wen_50 ? _GEN_7301 : data_5_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7334 = wen_50 ? _GEN_7302 : data_6_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7335 = wen_50 ? _GEN_7303 : data_7_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7336 = wen_50 ? _GEN_7304 : data_8_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7337 = wen_50 ? _GEN_7305 : data_9_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7338 = wen_50 ? _GEN_7306 : data_10_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7339 = wen_50 ? _GEN_7307 : data_11_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7340 = wen_50 ? _GEN_7308 : data_12_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7341 = wen_50 ? _GEN_7309 : data_13_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7342 = wen_50 ? _GEN_7310 : data_14_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7343 = wen_50 ? _GEN_7311 : data_15_6_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7344 = wen_50 ? _GEN_7312 : _GEN_3872; // @[Sbuffer.scala 160:18]
  wire  _GEN_7345 = wen_50 ? _GEN_7313 : _GEN_3873; // @[Sbuffer.scala 160:18]
  wire  _GEN_7346 = wen_50 ? _GEN_7314 : _GEN_3874; // @[Sbuffer.scala 160:18]
  wire  _GEN_7347 = wen_50 ? _GEN_7315 : _GEN_3875; // @[Sbuffer.scala 160:18]
  wire  _GEN_7348 = wen_50 ? _GEN_7316 : _GEN_3876; // @[Sbuffer.scala 160:18]
  wire  _GEN_7349 = wen_50 ? _GEN_7317 : _GEN_3877; // @[Sbuffer.scala 160:18]
  wire  _GEN_7350 = wen_50 ? _GEN_7318 : _GEN_3878; // @[Sbuffer.scala 160:18]
  wire  _GEN_7351 = wen_50 ? _GEN_7319 : _GEN_3879; // @[Sbuffer.scala 160:18]
  wire  _GEN_7352 = wen_50 ? _GEN_7320 : _GEN_3880; // @[Sbuffer.scala 160:18]
  wire  _GEN_7353 = wen_50 ? _GEN_7321 : _GEN_3881; // @[Sbuffer.scala 160:18]
  wire  _GEN_7354 = wen_50 ? _GEN_7322 : _GEN_3882; // @[Sbuffer.scala 160:18]
  wire  _GEN_7355 = wen_50 ? _GEN_7323 : _GEN_3883; // @[Sbuffer.scala 160:18]
  wire  _GEN_7356 = wen_50 ? _GEN_7324 : _GEN_3884; // @[Sbuffer.scala 160:18]
  wire  _GEN_7357 = wen_50 ? _GEN_7325 : _GEN_3885; // @[Sbuffer.scala 160:18]
  wire  _GEN_7358 = wen_50 ? _GEN_7326 : _GEN_3886; // @[Sbuffer.scala 160:18]
  wire  _GEN_7359 = wen_50 ? _GEN_7327 : _GEN_3887; // @[Sbuffer.scala 160:18]
  wire  _wen_T_207 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_51 = w_valid_s1_0 & _wen_T_207; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7360 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7361 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7362 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7363 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7364 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7365 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7366 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7367 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7368 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7369 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7370 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7371 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7372 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7373 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7374 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7375 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_6_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7376 = 4'h0 == w_addr_s1_0 | _GEN_3888; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7377 = 4'h1 == w_addr_s1_0 | _GEN_3889; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7378 = 4'h2 == w_addr_s1_0 | _GEN_3890; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7379 = 4'h3 == w_addr_s1_0 | _GEN_3891; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7380 = 4'h4 == w_addr_s1_0 | _GEN_3892; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7381 = 4'h5 == w_addr_s1_0 | _GEN_3893; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7382 = 4'h6 == w_addr_s1_0 | _GEN_3894; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7383 = 4'h7 == w_addr_s1_0 | _GEN_3895; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7384 = 4'h8 == w_addr_s1_0 | _GEN_3896; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7385 = 4'h9 == w_addr_s1_0 | _GEN_3897; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7386 = 4'ha == w_addr_s1_0 | _GEN_3898; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7387 = 4'hb == w_addr_s1_0 | _GEN_3899; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7388 = 4'hc == w_addr_s1_0 | _GEN_3900; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7389 = 4'hd == w_addr_s1_0 | _GEN_3901; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7390 = 4'he == w_addr_s1_0 | _GEN_3902; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7391 = 4'hf == w_addr_s1_0 | _GEN_3903; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7392 = wen_51 ? _GEN_7360 : data_0_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7393 = wen_51 ? _GEN_7361 : data_1_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7394 = wen_51 ? _GEN_7362 : data_2_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7395 = wen_51 ? _GEN_7363 : data_3_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7396 = wen_51 ? _GEN_7364 : data_4_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7397 = wen_51 ? _GEN_7365 : data_5_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7398 = wen_51 ? _GEN_7366 : data_6_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7399 = wen_51 ? _GEN_7367 : data_7_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7400 = wen_51 ? _GEN_7368 : data_8_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7401 = wen_51 ? _GEN_7369 : data_9_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7402 = wen_51 ? _GEN_7370 : data_10_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7403 = wen_51 ? _GEN_7371 : data_11_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7404 = wen_51 ? _GEN_7372 : data_12_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7405 = wen_51 ? _GEN_7373 : data_13_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7406 = wen_51 ? _GEN_7374 : data_14_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7407 = wen_51 ? _GEN_7375 : data_15_6_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7408 = wen_51 ? _GEN_7376 : _GEN_3888; // @[Sbuffer.scala 160:18]
  wire  _GEN_7409 = wen_51 ? _GEN_7377 : _GEN_3889; // @[Sbuffer.scala 160:18]
  wire  _GEN_7410 = wen_51 ? _GEN_7378 : _GEN_3890; // @[Sbuffer.scala 160:18]
  wire  _GEN_7411 = wen_51 ? _GEN_7379 : _GEN_3891; // @[Sbuffer.scala 160:18]
  wire  _GEN_7412 = wen_51 ? _GEN_7380 : _GEN_3892; // @[Sbuffer.scala 160:18]
  wire  _GEN_7413 = wen_51 ? _GEN_7381 : _GEN_3893; // @[Sbuffer.scala 160:18]
  wire  _GEN_7414 = wen_51 ? _GEN_7382 : _GEN_3894; // @[Sbuffer.scala 160:18]
  wire  _GEN_7415 = wen_51 ? _GEN_7383 : _GEN_3895; // @[Sbuffer.scala 160:18]
  wire  _GEN_7416 = wen_51 ? _GEN_7384 : _GEN_3896; // @[Sbuffer.scala 160:18]
  wire  _GEN_7417 = wen_51 ? _GEN_7385 : _GEN_3897; // @[Sbuffer.scala 160:18]
  wire  _GEN_7418 = wen_51 ? _GEN_7386 : _GEN_3898; // @[Sbuffer.scala 160:18]
  wire  _GEN_7419 = wen_51 ? _GEN_7387 : _GEN_3899; // @[Sbuffer.scala 160:18]
  wire  _GEN_7420 = wen_51 ? _GEN_7388 : _GEN_3900; // @[Sbuffer.scala 160:18]
  wire  _GEN_7421 = wen_51 ? _GEN_7389 : _GEN_3901; // @[Sbuffer.scala 160:18]
  wire  _GEN_7422 = wen_51 ? _GEN_7390 : _GEN_3902; // @[Sbuffer.scala 160:18]
  wire  _GEN_7423 = wen_51 ? _GEN_7391 : _GEN_3903; // @[Sbuffer.scala 160:18]
  wire  _wen_T_211 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_52 = w_valid_s1_0 & _wen_T_211; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7424 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7425 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7426 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7427 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7428 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7429 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7430 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7431 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7432 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7433 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7434 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7435 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7436 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7437 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7438 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7439 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_6_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7440 = 4'h0 == w_addr_s1_0 | _GEN_3904; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7441 = 4'h1 == w_addr_s1_0 | _GEN_3905; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7442 = 4'h2 == w_addr_s1_0 | _GEN_3906; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7443 = 4'h3 == w_addr_s1_0 | _GEN_3907; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7444 = 4'h4 == w_addr_s1_0 | _GEN_3908; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7445 = 4'h5 == w_addr_s1_0 | _GEN_3909; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7446 = 4'h6 == w_addr_s1_0 | _GEN_3910; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7447 = 4'h7 == w_addr_s1_0 | _GEN_3911; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7448 = 4'h8 == w_addr_s1_0 | _GEN_3912; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7449 = 4'h9 == w_addr_s1_0 | _GEN_3913; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7450 = 4'ha == w_addr_s1_0 | _GEN_3914; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7451 = 4'hb == w_addr_s1_0 | _GEN_3915; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7452 = 4'hc == w_addr_s1_0 | _GEN_3916; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7453 = 4'hd == w_addr_s1_0 | _GEN_3917; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7454 = 4'he == w_addr_s1_0 | _GEN_3918; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7455 = 4'hf == w_addr_s1_0 | _GEN_3919; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7456 = wen_52 ? _GEN_7424 : data_0_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7457 = wen_52 ? _GEN_7425 : data_1_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7458 = wen_52 ? _GEN_7426 : data_2_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7459 = wen_52 ? _GEN_7427 : data_3_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7460 = wen_52 ? _GEN_7428 : data_4_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7461 = wen_52 ? _GEN_7429 : data_5_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7462 = wen_52 ? _GEN_7430 : data_6_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7463 = wen_52 ? _GEN_7431 : data_7_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7464 = wen_52 ? _GEN_7432 : data_8_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7465 = wen_52 ? _GEN_7433 : data_9_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7466 = wen_52 ? _GEN_7434 : data_10_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7467 = wen_52 ? _GEN_7435 : data_11_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7468 = wen_52 ? _GEN_7436 : data_12_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7469 = wen_52 ? _GEN_7437 : data_13_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7470 = wen_52 ? _GEN_7438 : data_14_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7471 = wen_52 ? _GEN_7439 : data_15_6_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7472 = wen_52 ? _GEN_7440 : _GEN_3904; // @[Sbuffer.scala 160:18]
  wire  _GEN_7473 = wen_52 ? _GEN_7441 : _GEN_3905; // @[Sbuffer.scala 160:18]
  wire  _GEN_7474 = wen_52 ? _GEN_7442 : _GEN_3906; // @[Sbuffer.scala 160:18]
  wire  _GEN_7475 = wen_52 ? _GEN_7443 : _GEN_3907; // @[Sbuffer.scala 160:18]
  wire  _GEN_7476 = wen_52 ? _GEN_7444 : _GEN_3908; // @[Sbuffer.scala 160:18]
  wire  _GEN_7477 = wen_52 ? _GEN_7445 : _GEN_3909; // @[Sbuffer.scala 160:18]
  wire  _GEN_7478 = wen_52 ? _GEN_7446 : _GEN_3910; // @[Sbuffer.scala 160:18]
  wire  _GEN_7479 = wen_52 ? _GEN_7447 : _GEN_3911; // @[Sbuffer.scala 160:18]
  wire  _GEN_7480 = wen_52 ? _GEN_7448 : _GEN_3912; // @[Sbuffer.scala 160:18]
  wire  _GEN_7481 = wen_52 ? _GEN_7449 : _GEN_3913; // @[Sbuffer.scala 160:18]
  wire  _GEN_7482 = wen_52 ? _GEN_7450 : _GEN_3914; // @[Sbuffer.scala 160:18]
  wire  _GEN_7483 = wen_52 ? _GEN_7451 : _GEN_3915; // @[Sbuffer.scala 160:18]
  wire  _GEN_7484 = wen_52 ? _GEN_7452 : _GEN_3916; // @[Sbuffer.scala 160:18]
  wire  _GEN_7485 = wen_52 ? _GEN_7453 : _GEN_3917; // @[Sbuffer.scala 160:18]
  wire  _GEN_7486 = wen_52 ? _GEN_7454 : _GEN_3918; // @[Sbuffer.scala 160:18]
  wire  _GEN_7487 = wen_52 ? _GEN_7455 : _GEN_3919; // @[Sbuffer.scala 160:18]
  wire  _wen_T_215 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_53 = w_valid_s1_0 & _wen_T_215; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7488 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7489 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7490 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7491 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7492 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7493 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7494 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7495 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7496 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7497 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7498 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7499 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7500 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7501 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7502 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7503 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_6_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7504 = 4'h0 == w_addr_s1_0 | _GEN_3920; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7505 = 4'h1 == w_addr_s1_0 | _GEN_3921; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7506 = 4'h2 == w_addr_s1_0 | _GEN_3922; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7507 = 4'h3 == w_addr_s1_0 | _GEN_3923; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7508 = 4'h4 == w_addr_s1_0 | _GEN_3924; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7509 = 4'h5 == w_addr_s1_0 | _GEN_3925; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7510 = 4'h6 == w_addr_s1_0 | _GEN_3926; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7511 = 4'h7 == w_addr_s1_0 | _GEN_3927; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7512 = 4'h8 == w_addr_s1_0 | _GEN_3928; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7513 = 4'h9 == w_addr_s1_0 | _GEN_3929; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7514 = 4'ha == w_addr_s1_0 | _GEN_3930; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7515 = 4'hb == w_addr_s1_0 | _GEN_3931; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7516 = 4'hc == w_addr_s1_0 | _GEN_3932; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7517 = 4'hd == w_addr_s1_0 | _GEN_3933; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7518 = 4'he == w_addr_s1_0 | _GEN_3934; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7519 = 4'hf == w_addr_s1_0 | _GEN_3935; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7520 = wen_53 ? _GEN_7488 : data_0_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7521 = wen_53 ? _GEN_7489 : data_1_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7522 = wen_53 ? _GEN_7490 : data_2_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7523 = wen_53 ? _GEN_7491 : data_3_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7524 = wen_53 ? _GEN_7492 : data_4_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7525 = wen_53 ? _GEN_7493 : data_5_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7526 = wen_53 ? _GEN_7494 : data_6_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7527 = wen_53 ? _GEN_7495 : data_7_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7528 = wen_53 ? _GEN_7496 : data_8_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7529 = wen_53 ? _GEN_7497 : data_9_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7530 = wen_53 ? _GEN_7498 : data_10_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7531 = wen_53 ? _GEN_7499 : data_11_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7532 = wen_53 ? _GEN_7500 : data_12_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7533 = wen_53 ? _GEN_7501 : data_13_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7534 = wen_53 ? _GEN_7502 : data_14_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7535 = wen_53 ? _GEN_7503 : data_15_6_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7536 = wen_53 ? _GEN_7504 : _GEN_3920; // @[Sbuffer.scala 160:18]
  wire  _GEN_7537 = wen_53 ? _GEN_7505 : _GEN_3921; // @[Sbuffer.scala 160:18]
  wire  _GEN_7538 = wen_53 ? _GEN_7506 : _GEN_3922; // @[Sbuffer.scala 160:18]
  wire  _GEN_7539 = wen_53 ? _GEN_7507 : _GEN_3923; // @[Sbuffer.scala 160:18]
  wire  _GEN_7540 = wen_53 ? _GEN_7508 : _GEN_3924; // @[Sbuffer.scala 160:18]
  wire  _GEN_7541 = wen_53 ? _GEN_7509 : _GEN_3925; // @[Sbuffer.scala 160:18]
  wire  _GEN_7542 = wen_53 ? _GEN_7510 : _GEN_3926; // @[Sbuffer.scala 160:18]
  wire  _GEN_7543 = wen_53 ? _GEN_7511 : _GEN_3927; // @[Sbuffer.scala 160:18]
  wire  _GEN_7544 = wen_53 ? _GEN_7512 : _GEN_3928; // @[Sbuffer.scala 160:18]
  wire  _GEN_7545 = wen_53 ? _GEN_7513 : _GEN_3929; // @[Sbuffer.scala 160:18]
  wire  _GEN_7546 = wen_53 ? _GEN_7514 : _GEN_3930; // @[Sbuffer.scala 160:18]
  wire  _GEN_7547 = wen_53 ? _GEN_7515 : _GEN_3931; // @[Sbuffer.scala 160:18]
  wire  _GEN_7548 = wen_53 ? _GEN_7516 : _GEN_3932; // @[Sbuffer.scala 160:18]
  wire  _GEN_7549 = wen_53 ? _GEN_7517 : _GEN_3933; // @[Sbuffer.scala 160:18]
  wire  _GEN_7550 = wen_53 ? _GEN_7518 : _GEN_3934; // @[Sbuffer.scala 160:18]
  wire  _GEN_7551 = wen_53 ? _GEN_7519 : _GEN_3935; // @[Sbuffer.scala 160:18]
  wire  _wen_T_219 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_54 = w_valid_s1_0 & _wen_T_219; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7552 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7553 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7554 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7555 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7556 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7557 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7558 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7559 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7560 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7561 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7562 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7563 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7564 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7565 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7566 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7567 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_6_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7568 = 4'h0 == w_addr_s1_0 | _GEN_3936; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7569 = 4'h1 == w_addr_s1_0 | _GEN_3937; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7570 = 4'h2 == w_addr_s1_0 | _GEN_3938; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7571 = 4'h3 == w_addr_s1_0 | _GEN_3939; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7572 = 4'h4 == w_addr_s1_0 | _GEN_3940; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7573 = 4'h5 == w_addr_s1_0 | _GEN_3941; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7574 = 4'h6 == w_addr_s1_0 | _GEN_3942; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7575 = 4'h7 == w_addr_s1_0 | _GEN_3943; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7576 = 4'h8 == w_addr_s1_0 | _GEN_3944; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7577 = 4'h9 == w_addr_s1_0 | _GEN_3945; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7578 = 4'ha == w_addr_s1_0 | _GEN_3946; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7579 = 4'hb == w_addr_s1_0 | _GEN_3947; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7580 = 4'hc == w_addr_s1_0 | _GEN_3948; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7581 = 4'hd == w_addr_s1_0 | _GEN_3949; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7582 = 4'he == w_addr_s1_0 | _GEN_3950; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7583 = 4'hf == w_addr_s1_0 | _GEN_3951; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7584 = wen_54 ? _GEN_7552 : data_0_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7585 = wen_54 ? _GEN_7553 : data_1_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7586 = wen_54 ? _GEN_7554 : data_2_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7587 = wen_54 ? _GEN_7555 : data_3_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7588 = wen_54 ? _GEN_7556 : data_4_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7589 = wen_54 ? _GEN_7557 : data_5_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7590 = wen_54 ? _GEN_7558 : data_6_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7591 = wen_54 ? _GEN_7559 : data_7_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7592 = wen_54 ? _GEN_7560 : data_8_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7593 = wen_54 ? _GEN_7561 : data_9_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7594 = wen_54 ? _GEN_7562 : data_10_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7595 = wen_54 ? _GEN_7563 : data_11_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7596 = wen_54 ? _GEN_7564 : data_12_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7597 = wen_54 ? _GEN_7565 : data_13_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7598 = wen_54 ? _GEN_7566 : data_14_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7599 = wen_54 ? _GEN_7567 : data_15_6_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7600 = wen_54 ? _GEN_7568 : _GEN_3936; // @[Sbuffer.scala 160:18]
  wire  _GEN_7601 = wen_54 ? _GEN_7569 : _GEN_3937; // @[Sbuffer.scala 160:18]
  wire  _GEN_7602 = wen_54 ? _GEN_7570 : _GEN_3938; // @[Sbuffer.scala 160:18]
  wire  _GEN_7603 = wen_54 ? _GEN_7571 : _GEN_3939; // @[Sbuffer.scala 160:18]
  wire  _GEN_7604 = wen_54 ? _GEN_7572 : _GEN_3940; // @[Sbuffer.scala 160:18]
  wire  _GEN_7605 = wen_54 ? _GEN_7573 : _GEN_3941; // @[Sbuffer.scala 160:18]
  wire  _GEN_7606 = wen_54 ? _GEN_7574 : _GEN_3942; // @[Sbuffer.scala 160:18]
  wire  _GEN_7607 = wen_54 ? _GEN_7575 : _GEN_3943; // @[Sbuffer.scala 160:18]
  wire  _GEN_7608 = wen_54 ? _GEN_7576 : _GEN_3944; // @[Sbuffer.scala 160:18]
  wire  _GEN_7609 = wen_54 ? _GEN_7577 : _GEN_3945; // @[Sbuffer.scala 160:18]
  wire  _GEN_7610 = wen_54 ? _GEN_7578 : _GEN_3946; // @[Sbuffer.scala 160:18]
  wire  _GEN_7611 = wen_54 ? _GEN_7579 : _GEN_3947; // @[Sbuffer.scala 160:18]
  wire  _GEN_7612 = wen_54 ? _GEN_7580 : _GEN_3948; // @[Sbuffer.scala 160:18]
  wire  _GEN_7613 = wen_54 ? _GEN_7581 : _GEN_3949; // @[Sbuffer.scala 160:18]
  wire  _GEN_7614 = wen_54 ? _GEN_7582 : _GEN_3950; // @[Sbuffer.scala 160:18]
  wire  _GEN_7615 = wen_54 ? _GEN_7583 : _GEN_3951; // @[Sbuffer.scala 160:18]
  wire  _wen_T_223 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h6 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_55 = w_valid_s1_0 & _wen_T_223; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7616 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7617 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7618 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7619 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7620 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7621 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7622 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7623 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7624 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7625 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7626 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7627 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7628 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7629 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7630 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7631 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_6_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7632 = 4'h0 == w_addr_s1_0 | _GEN_3952; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7633 = 4'h1 == w_addr_s1_0 | _GEN_3953; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7634 = 4'h2 == w_addr_s1_0 | _GEN_3954; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7635 = 4'h3 == w_addr_s1_0 | _GEN_3955; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7636 = 4'h4 == w_addr_s1_0 | _GEN_3956; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7637 = 4'h5 == w_addr_s1_0 | _GEN_3957; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7638 = 4'h6 == w_addr_s1_0 | _GEN_3958; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7639 = 4'h7 == w_addr_s1_0 | _GEN_3959; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7640 = 4'h8 == w_addr_s1_0 | _GEN_3960; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7641 = 4'h9 == w_addr_s1_0 | _GEN_3961; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7642 = 4'ha == w_addr_s1_0 | _GEN_3962; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7643 = 4'hb == w_addr_s1_0 | _GEN_3963; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7644 = 4'hc == w_addr_s1_0 | _GEN_3964; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7645 = 4'hd == w_addr_s1_0 | _GEN_3965; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7646 = 4'he == w_addr_s1_0 | _GEN_3966; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7647 = 4'hf == w_addr_s1_0 | _GEN_3967; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7648 = wen_55 ? _GEN_7616 : data_0_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7649 = wen_55 ? _GEN_7617 : data_1_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7650 = wen_55 ? _GEN_7618 : data_2_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7651 = wen_55 ? _GEN_7619 : data_3_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7652 = wen_55 ? _GEN_7620 : data_4_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7653 = wen_55 ? _GEN_7621 : data_5_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7654 = wen_55 ? _GEN_7622 : data_6_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7655 = wen_55 ? _GEN_7623 : data_7_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7656 = wen_55 ? _GEN_7624 : data_8_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7657 = wen_55 ? _GEN_7625 : data_9_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7658 = wen_55 ? _GEN_7626 : data_10_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7659 = wen_55 ? _GEN_7627 : data_11_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7660 = wen_55 ? _GEN_7628 : data_12_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7661 = wen_55 ? _GEN_7629 : data_13_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7662 = wen_55 ? _GEN_7630 : data_14_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7663 = wen_55 ? _GEN_7631 : data_15_6_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7664 = wen_55 ? _GEN_7632 : _GEN_3952; // @[Sbuffer.scala 160:18]
  wire  _GEN_7665 = wen_55 ? _GEN_7633 : _GEN_3953; // @[Sbuffer.scala 160:18]
  wire  _GEN_7666 = wen_55 ? _GEN_7634 : _GEN_3954; // @[Sbuffer.scala 160:18]
  wire  _GEN_7667 = wen_55 ? _GEN_7635 : _GEN_3955; // @[Sbuffer.scala 160:18]
  wire  _GEN_7668 = wen_55 ? _GEN_7636 : _GEN_3956; // @[Sbuffer.scala 160:18]
  wire  _GEN_7669 = wen_55 ? _GEN_7637 : _GEN_3957; // @[Sbuffer.scala 160:18]
  wire  _GEN_7670 = wen_55 ? _GEN_7638 : _GEN_3958; // @[Sbuffer.scala 160:18]
  wire  _GEN_7671 = wen_55 ? _GEN_7639 : _GEN_3959; // @[Sbuffer.scala 160:18]
  wire  _GEN_7672 = wen_55 ? _GEN_7640 : _GEN_3960; // @[Sbuffer.scala 160:18]
  wire  _GEN_7673 = wen_55 ? _GEN_7641 : _GEN_3961; // @[Sbuffer.scala 160:18]
  wire  _GEN_7674 = wen_55 ? _GEN_7642 : _GEN_3962; // @[Sbuffer.scala 160:18]
  wire  _GEN_7675 = wen_55 ? _GEN_7643 : _GEN_3963; // @[Sbuffer.scala 160:18]
  wire  _GEN_7676 = wen_55 ? _GEN_7644 : _GEN_3964; // @[Sbuffer.scala 160:18]
  wire  _GEN_7677 = wen_55 ? _GEN_7645 : _GEN_3965; // @[Sbuffer.scala 160:18]
  wire  _GEN_7678 = wen_55 ? _GEN_7646 : _GEN_3966; // @[Sbuffer.scala 160:18]
  wire  _GEN_7679 = wen_55 ? _GEN_7647 : _GEN_3967; // @[Sbuffer.scala 160:18]
  wire  _wen_T_227 = w_mask_s1_0[0] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_56 = w_valid_s1_0 & _wen_T_227; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7680 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_0_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7681 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_1_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7682 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_2_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7683 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_3_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7684 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_4_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7685 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_5_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7686 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_6_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7687 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_7_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7688 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_8_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7689 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[7:0] : data_9_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7690 = 4'ha == w_addr_s1_0 ? w_data_s1_0[7:0] : data_10_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7691 = 4'hb == w_addr_s1_0 ? w_data_s1_0[7:0] : data_11_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7692 = 4'hc == w_addr_s1_0 ? w_data_s1_0[7:0] : data_12_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7693 = 4'hd == w_addr_s1_0 ? w_data_s1_0[7:0] : data_13_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7694 = 4'he == w_addr_s1_0 ? w_data_s1_0[7:0] : data_14_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7695 = 4'hf == w_addr_s1_0 ? w_data_s1_0[7:0] : data_15_7_0; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7696 = 4'h0 == w_addr_s1_0 | _GEN_3968; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7697 = 4'h1 == w_addr_s1_0 | _GEN_3969; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7698 = 4'h2 == w_addr_s1_0 | _GEN_3970; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7699 = 4'h3 == w_addr_s1_0 | _GEN_3971; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7700 = 4'h4 == w_addr_s1_0 | _GEN_3972; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7701 = 4'h5 == w_addr_s1_0 | _GEN_3973; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7702 = 4'h6 == w_addr_s1_0 | _GEN_3974; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7703 = 4'h7 == w_addr_s1_0 | _GEN_3975; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7704 = 4'h8 == w_addr_s1_0 | _GEN_3976; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7705 = 4'h9 == w_addr_s1_0 | _GEN_3977; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7706 = 4'ha == w_addr_s1_0 | _GEN_3978; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7707 = 4'hb == w_addr_s1_0 | _GEN_3979; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7708 = 4'hc == w_addr_s1_0 | _GEN_3980; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7709 = 4'hd == w_addr_s1_0 | _GEN_3981; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7710 = 4'he == w_addr_s1_0 | _GEN_3982; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7711 = 4'hf == w_addr_s1_0 | _GEN_3983; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7712 = wen_56 ? _GEN_7680 : data_0_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7713 = wen_56 ? _GEN_7681 : data_1_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7714 = wen_56 ? _GEN_7682 : data_2_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7715 = wen_56 ? _GEN_7683 : data_3_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7716 = wen_56 ? _GEN_7684 : data_4_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7717 = wen_56 ? _GEN_7685 : data_5_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7718 = wen_56 ? _GEN_7686 : data_6_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7719 = wen_56 ? _GEN_7687 : data_7_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7720 = wen_56 ? _GEN_7688 : data_8_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7721 = wen_56 ? _GEN_7689 : data_9_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7722 = wen_56 ? _GEN_7690 : data_10_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7723 = wen_56 ? _GEN_7691 : data_11_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7724 = wen_56 ? _GEN_7692 : data_12_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7725 = wen_56 ? _GEN_7693 : data_13_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7726 = wen_56 ? _GEN_7694 : data_14_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7727 = wen_56 ? _GEN_7695 : data_15_7_0; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7728 = wen_56 ? _GEN_7696 : _GEN_3968; // @[Sbuffer.scala 160:18]
  wire  _GEN_7729 = wen_56 ? _GEN_7697 : _GEN_3969; // @[Sbuffer.scala 160:18]
  wire  _GEN_7730 = wen_56 ? _GEN_7698 : _GEN_3970; // @[Sbuffer.scala 160:18]
  wire  _GEN_7731 = wen_56 ? _GEN_7699 : _GEN_3971; // @[Sbuffer.scala 160:18]
  wire  _GEN_7732 = wen_56 ? _GEN_7700 : _GEN_3972; // @[Sbuffer.scala 160:18]
  wire  _GEN_7733 = wen_56 ? _GEN_7701 : _GEN_3973; // @[Sbuffer.scala 160:18]
  wire  _GEN_7734 = wen_56 ? _GEN_7702 : _GEN_3974; // @[Sbuffer.scala 160:18]
  wire  _GEN_7735 = wen_56 ? _GEN_7703 : _GEN_3975; // @[Sbuffer.scala 160:18]
  wire  _GEN_7736 = wen_56 ? _GEN_7704 : _GEN_3976; // @[Sbuffer.scala 160:18]
  wire  _GEN_7737 = wen_56 ? _GEN_7705 : _GEN_3977; // @[Sbuffer.scala 160:18]
  wire  _GEN_7738 = wen_56 ? _GEN_7706 : _GEN_3978; // @[Sbuffer.scala 160:18]
  wire  _GEN_7739 = wen_56 ? _GEN_7707 : _GEN_3979; // @[Sbuffer.scala 160:18]
  wire  _GEN_7740 = wen_56 ? _GEN_7708 : _GEN_3980; // @[Sbuffer.scala 160:18]
  wire  _GEN_7741 = wen_56 ? _GEN_7709 : _GEN_3981; // @[Sbuffer.scala 160:18]
  wire  _GEN_7742 = wen_56 ? _GEN_7710 : _GEN_3982; // @[Sbuffer.scala 160:18]
  wire  _GEN_7743 = wen_56 ? _GEN_7711 : _GEN_3983; // @[Sbuffer.scala 160:18]
  wire  _wen_T_231 = w_mask_s1_0[1] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_57 = w_valid_s1_0 & _wen_T_231; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7744 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_0_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7745 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_1_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7746 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_2_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7747 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_3_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7748 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_4_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7749 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_5_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7750 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_6_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7751 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_7_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7752 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_8_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7753 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[15:8] : data_9_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7754 = 4'ha == w_addr_s1_0 ? w_data_s1_0[15:8] : data_10_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7755 = 4'hb == w_addr_s1_0 ? w_data_s1_0[15:8] : data_11_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7756 = 4'hc == w_addr_s1_0 ? w_data_s1_0[15:8] : data_12_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7757 = 4'hd == w_addr_s1_0 ? w_data_s1_0[15:8] : data_13_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7758 = 4'he == w_addr_s1_0 ? w_data_s1_0[15:8] : data_14_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7759 = 4'hf == w_addr_s1_0 ? w_data_s1_0[15:8] : data_15_7_1; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7760 = 4'h0 == w_addr_s1_0 | _GEN_3984; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7761 = 4'h1 == w_addr_s1_0 | _GEN_3985; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7762 = 4'h2 == w_addr_s1_0 | _GEN_3986; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7763 = 4'h3 == w_addr_s1_0 | _GEN_3987; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7764 = 4'h4 == w_addr_s1_0 | _GEN_3988; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7765 = 4'h5 == w_addr_s1_0 | _GEN_3989; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7766 = 4'h6 == w_addr_s1_0 | _GEN_3990; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7767 = 4'h7 == w_addr_s1_0 | _GEN_3991; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7768 = 4'h8 == w_addr_s1_0 | _GEN_3992; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7769 = 4'h9 == w_addr_s1_0 | _GEN_3993; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7770 = 4'ha == w_addr_s1_0 | _GEN_3994; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7771 = 4'hb == w_addr_s1_0 | _GEN_3995; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7772 = 4'hc == w_addr_s1_0 | _GEN_3996; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7773 = 4'hd == w_addr_s1_0 | _GEN_3997; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7774 = 4'he == w_addr_s1_0 | _GEN_3998; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7775 = 4'hf == w_addr_s1_0 | _GEN_3999; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7776 = wen_57 ? _GEN_7744 : data_0_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7777 = wen_57 ? _GEN_7745 : data_1_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7778 = wen_57 ? _GEN_7746 : data_2_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7779 = wen_57 ? _GEN_7747 : data_3_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7780 = wen_57 ? _GEN_7748 : data_4_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7781 = wen_57 ? _GEN_7749 : data_5_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7782 = wen_57 ? _GEN_7750 : data_6_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7783 = wen_57 ? _GEN_7751 : data_7_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7784 = wen_57 ? _GEN_7752 : data_8_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7785 = wen_57 ? _GEN_7753 : data_9_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7786 = wen_57 ? _GEN_7754 : data_10_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7787 = wen_57 ? _GEN_7755 : data_11_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7788 = wen_57 ? _GEN_7756 : data_12_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7789 = wen_57 ? _GEN_7757 : data_13_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7790 = wen_57 ? _GEN_7758 : data_14_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7791 = wen_57 ? _GEN_7759 : data_15_7_1; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7792 = wen_57 ? _GEN_7760 : _GEN_3984; // @[Sbuffer.scala 160:18]
  wire  _GEN_7793 = wen_57 ? _GEN_7761 : _GEN_3985; // @[Sbuffer.scala 160:18]
  wire  _GEN_7794 = wen_57 ? _GEN_7762 : _GEN_3986; // @[Sbuffer.scala 160:18]
  wire  _GEN_7795 = wen_57 ? _GEN_7763 : _GEN_3987; // @[Sbuffer.scala 160:18]
  wire  _GEN_7796 = wen_57 ? _GEN_7764 : _GEN_3988; // @[Sbuffer.scala 160:18]
  wire  _GEN_7797 = wen_57 ? _GEN_7765 : _GEN_3989; // @[Sbuffer.scala 160:18]
  wire  _GEN_7798 = wen_57 ? _GEN_7766 : _GEN_3990; // @[Sbuffer.scala 160:18]
  wire  _GEN_7799 = wen_57 ? _GEN_7767 : _GEN_3991; // @[Sbuffer.scala 160:18]
  wire  _GEN_7800 = wen_57 ? _GEN_7768 : _GEN_3992; // @[Sbuffer.scala 160:18]
  wire  _GEN_7801 = wen_57 ? _GEN_7769 : _GEN_3993; // @[Sbuffer.scala 160:18]
  wire  _GEN_7802 = wen_57 ? _GEN_7770 : _GEN_3994; // @[Sbuffer.scala 160:18]
  wire  _GEN_7803 = wen_57 ? _GEN_7771 : _GEN_3995; // @[Sbuffer.scala 160:18]
  wire  _GEN_7804 = wen_57 ? _GEN_7772 : _GEN_3996; // @[Sbuffer.scala 160:18]
  wire  _GEN_7805 = wen_57 ? _GEN_7773 : _GEN_3997; // @[Sbuffer.scala 160:18]
  wire  _GEN_7806 = wen_57 ? _GEN_7774 : _GEN_3998; // @[Sbuffer.scala 160:18]
  wire  _GEN_7807 = wen_57 ? _GEN_7775 : _GEN_3999; // @[Sbuffer.scala 160:18]
  wire  _wen_T_235 = w_mask_s1_0[2] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_58 = w_valid_s1_0 & _wen_T_235; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7808 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_0_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7809 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_1_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7810 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_2_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7811 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_3_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7812 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_4_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7813 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_5_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7814 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_6_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7815 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_7_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7816 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_8_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7817 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[23:16] : data_9_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7818 = 4'ha == w_addr_s1_0 ? w_data_s1_0[23:16] : data_10_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7819 = 4'hb == w_addr_s1_0 ? w_data_s1_0[23:16] : data_11_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7820 = 4'hc == w_addr_s1_0 ? w_data_s1_0[23:16] : data_12_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7821 = 4'hd == w_addr_s1_0 ? w_data_s1_0[23:16] : data_13_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7822 = 4'he == w_addr_s1_0 ? w_data_s1_0[23:16] : data_14_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7823 = 4'hf == w_addr_s1_0 ? w_data_s1_0[23:16] : data_15_7_2; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7824 = 4'h0 == w_addr_s1_0 | _GEN_4000; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7825 = 4'h1 == w_addr_s1_0 | _GEN_4001; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7826 = 4'h2 == w_addr_s1_0 | _GEN_4002; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7827 = 4'h3 == w_addr_s1_0 | _GEN_4003; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7828 = 4'h4 == w_addr_s1_0 | _GEN_4004; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7829 = 4'h5 == w_addr_s1_0 | _GEN_4005; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7830 = 4'h6 == w_addr_s1_0 | _GEN_4006; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7831 = 4'h7 == w_addr_s1_0 | _GEN_4007; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7832 = 4'h8 == w_addr_s1_0 | _GEN_4008; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7833 = 4'h9 == w_addr_s1_0 | _GEN_4009; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7834 = 4'ha == w_addr_s1_0 | _GEN_4010; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7835 = 4'hb == w_addr_s1_0 | _GEN_4011; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7836 = 4'hc == w_addr_s1_0 | _GEN_4012; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7837 = 4'hd == w_addr_s1_0 | _GEN_4013; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7838 = 4'he == w_addr_s1_0 | _GEN_4014; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7839 = 4'hf == w_addr_s1_0 | _GEN_4015; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7840 = wen_58 ? _GEN_7808 : data_0_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7841 = wen_58 ? _GEN_7809 : data_1_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7842 = wen_58 ? _GEN_7810 : data_2_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7843 = wen_58 ? _GEN_7811 : data_3_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7844 = wen_58 ? _GEN_7812 : data_4_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7845 = wen_58 ? _GEN_7813 : data_5_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7846 = wen_58 ? _GEN_7814 : data_6_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7847 = wen_58 ? _GEN_7815 : data_7_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7848 = wen_58 ? _GEN_7816 : data_8_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7849 = wen_58 ? _GEN_7817 : data_9_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7850 = wen_58 ? _GEN_7818 : data_10_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7851 = wen_58 ? _GEN_7819 : data_11_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7852 = wen_58 ? _GEN_7820 : data_12_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7853 = wen_58 ? _GEN_7821 : data_13_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7854 = wen_58 ? _GEN_7822 : data_14_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7855 = wen_58 ? _GEN_7823 : data_15_7_2; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7856 = wen_58 ? _GEN_7824 : _GEN_4000; // @[Sbuffer.scala 160:18]
  wire  _GEN_7857 = wen_58 ? _GEN_7825 : _GEN_4001; // @[Sbuffer.scala 160:18]
  wire  _GEN_7858 = wen_58 ? _GEN_7826 : _GEN_4002; // @[Sbuffer.scala 160:18]
  wire  _GEN_7859 = wen_58 ? _GEN_7827 : _GEN_4003; // @[Sbuffer.scala 160:18]
  wire  _GEN_7860 = wen_58 ? _GEN_7828 : _GEN_4004; // @[Sbuffer.scala 160:18]
  wire  _GEN_7861 = wen_58 ? _GEN_7829 : _GEN_4005; // @[Sbuffer.scala 160:18]
  wire  _GEN_7862 = wen_58 ? _GEN_7830 : _GEN_4006; // @[Sbuffer.scala 160:18]
  wire  _GEN_7863 = wen_58 ? _GEN_7831 : _GEN_4007; // @[Sbuffer.scala 160:18]
  wire  _GEN_7864 = wen_58 ? _GEN_7832 : _GEN_4008; // @[Sbuffer.scala 160:18]
  wire  _GEN_7865 = wen_58 ? _GEN_7833 : _GEN_4009; // @[Sbuffer.scala 160:18]
  wire  _GEN_7866 = wen_58 ? _GEN_7834 : _GEN_4010; // @[Sbuffer.scala 160:18]
  wire  _GEN_7867 = wen_58 ? _GEN_7835 : _GEN_4011; // @[Sbuffer.scala 160:18]
  wire  _GEN_7868 = wen_58 ? _GEN_7836 : _GEN_4012; // @[Sbuffer.scala 160:18]
  wire  _GEN_7869 = wen_58 ? _GEN_7837 : _GEN_4013; // @[Sbuffer.scala 160:18]
  wire  _GEN_7870 = wen_58 ? _GEN_7838 : _GEN_4014; // @[Sbuffer.scala 160:18]
  wire  _GEN_7871 = wen_58 ? _GEN_7839 : _GEN_4015; // @[Sbuffer.scala 160:18]
  wire  _wen_T_239 = w_mask_s1_0[3] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_59 = w_valid_s1_0 & _wen_T_239; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7872 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_0_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7873 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_1_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7874 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_2_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7875 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_3_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7876 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_4_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7877 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_5_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7878 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_6_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7879 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_7_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7880 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_8_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7881 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[31:24] : data_9_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7882 = 4'ha == w_addr_s1_0 ? w_data_s1_0[31:24] : data_10_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7883 = 4'hb == w_addr_s1_0 ? w_data_s1_0[31:24] : data_11_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7884 = 4'hc == w_addr_s1_0 ? w_data_s1_0[31:24] : data_12_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7885 = 4'hd == w_addr_s1_0 ? w_data_s1_0[31:24] : data_13_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7886 = 4'he == w_addr_s1_0 ? w_data_s1_0[31:24] : data_14_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7887 = 4'hf == w_addr_s1_0 ? w_data_s1_0[31:24] : data_15_7_3; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7888 = 4'h0 == w_addr_s1_0 | _GEN_4016; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7889 = 4'h1 == w_addr_s1_0 | _GEN_4017; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7890 = 4'h2 == w_addr_s1_0 | _GEN_4018; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7891 = 4'h3 == w_addr_s1_0 | _GEN_4019; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7892 = 4'h4 == w_addr_s1_0 | _GEN_4020; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7893 = 4'h5 == w_addr_s1_0 | _GEN_4021; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7894 = 4'h6 == w_addr_s1_0 | _GEN_4022; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7895 = 4'h7 == w_addr_s1_0 | _GEN_4023; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7896 = 4'h8 == w_addr_s1_0 | _GEN_4024; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7897 = 4'h9 == w_addr_s1_0 | _GEN_4025; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7898 = 4'ha == w_addr_s1_0 | _GEN_4026; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7899 = 4'hb == w_addr_s1_0 | _GEN_4027; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7900 = 4'hc == w_addr_s1_0 | _GEN_4028; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7901 = 4'hd == w_addr_s1_0 | _GEN_4029; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7902 = 4'he == w_addr_s1_0 | _GEN_4030; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7903 = 4'hf == w_addr_s1_0 | _GEN_4031; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7904 = wen_59 ? _GEN_7872 : data_0_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7905 = wen_59 ? _GEN_7873 : data_1_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7906 = wen_59 ? _GEN_7874 : data_2_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7907 = wen_59 ? _GEN_7875 : data_3_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7908 = wen_59 ? _GEN_7876 : data_4_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7909 = wen_59 ? _GEN_7877 : data_5_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7910 = wen_59 ? _GEN_7878 : data_6_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7911 = wen_59 ? _GEN_7879 : data_7_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7912 = wen_59 ? _GEN_7880 : data_8_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7913 = wen_59 ? _GEN_7881 : data_9_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7914 = wen_59 ? _GEN_7882 : data_10_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7915 = wen_59 ? _GEN_7883 : data_11_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7916 = wen_59 ? _GEN_7884 : data_12_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7917 = wen_59 ? _GEN_7885 : data_13_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7918 = wen_59 ? _GEN_7886 : data_14_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7919 = wen_59 ? _GEN_7887 : data_15_7_3; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7920 = wen_59 ? _GEN_7888 : _GEN_4016; // @[Sbuffer.scala 160:18]
  wire  _GEN_7921 = wen_59 ? _GEN_7889 : _GEN_4017; // @[Sbuffer.scala 160:18]
  wire  _GEN_7922 = wen_59 ? _GEN_7890 : _GEN_4018; // @[Sbuffer.scala 160:18]
  wire  _GEN_7923 = wen_59 ? _GEN_7891 : _GEN_4019; // @[Sbuffer.scala 160:18]
  wire  _GEN_7924 = wen_59 ? _GEN_7892 : _GEN_4020; // @[Sbuffer.scala 160:18]
  wire  _GEN_7925 = wen_59 ? _GEN_7893 : _GEN_4021; // @[Sbuffer.scala 160:18]
  wire  _GEN_7926 = wen_59 ? _GEN_7894 : _GEN_4022; // @[Sbuffer.scala 160:18]
  wire  _GEN_7927 = wen_59 ? _GEN_7895 : _GEN_4023; // @[Sbuffer.scala 160:18]
  wire  _GEN_7928 = wen_59 ? _GEN_7896 : _GEN_4024; // @[Sbuffer.scala 160:18]
  wire  _GEN_7929 = wen_59 ? _GEN_7897 : _GEN_4025; // @[Sbuffer.scala 160:18]
  wire  _GEN_7930 = wen_59 ? _GEN_7898 : _GEN_4026; // @[Sbuffer.scala 160:18]
  wire  _GEN_7931 = wen_59 ? _GEN_7899 : _GEN_4027; // @[Sbuffer.scala 160:18]
  wire  _GEN_7932 = wen_59 ? _GEN_7900 : _GEN_4028; // @[Sbuffer.scala 160:18]
  wire  _GEN_7933 = wen_59 ? _GEN_7901 : _GEN_4029; // @[Sbuffer.scala 160:18]
  wire  _GEN_7934 = wen_59 ? _GEN_7902 : _GEN_4030; // @[Sbuffer.scala 160:18]
  wire  _GEN_7935 = wen_59 ? _GEN_7903 : _GEN_4031; // @[Sbuffer.scala 160:18]
  wire  _wen_T_243 = w_mask_s1_0[4] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_60 = w_valid_s1_0 & _wen_T_243; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_7936 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_0_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7937 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_1_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7938 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_2_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7939 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_3_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7940 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_4_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7941 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_5_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7942 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_6_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7943 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_7_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7944 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_8_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7945 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[39:32] : data_9_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7946 = 4'ha == w_addr_s1_0 ? w_data_s1_0[39:32] : data_10_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7947 = 4'hb == w_addr_s1_0 ? w_data_s1_0[39:32] : data_11_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7948 = 4'hc == w_addr_s1_0 ? w_data_s1_0[39:32] : data_12_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7949 = 4'hd == w_addr_s1_0 ? w_data_s1_0[39:32] : data_13_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7950 = 4'he == w_addr_s1_0 ? w_data_s1_0[39:32] : data_14_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_7951 = 4'hf == w_addr_s1_0 ? w_data_s1_0[39:32] : data_15_7_4; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_7952 = 4'h0 == w_addr_s1_0 | _GEN_4032; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7953 = 4'h1 == w_addr_s1_0 | _GEN_4033; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7954 = 4'h2 == w_addr_s1_0 | _GEN_4034; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7955 = 4'h3 == w_addr_s1_0 | _GEN_4035; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7956 = 4'h4 == w_addr_s1_0 | _GEN_4036; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7957 = 4'h5 == w_addr_s1_0 | _GEN_4037; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7958 = 4'h6 == w_addr_s1_0 | _GEN_4038; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7959 = 4'h7 == w_addr_s1_0 | _GEN_4039; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7960 = 4'h8 == w_addr_s1_0 | _GEN_4040; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7961 = 4'h9 == w_addr_s1_0 | _GEN_4041; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7962 = 4'ha == w_addr_s1_0 | _GEN_4042; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7963 = 4'hb == w_addr_s1_0 | _GEN_4043; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7964 = 4'hc == w_addr_s1_0 | _GEN_4044; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7965 = 4'hd == w_addr_s1_0 | _GEN_4045; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7966 = 4'he == w_addr_s1_0 | _GEN_4046; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_7967 = 4'hf == w_addr_s1_0 | _GEN_4047; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_7968 = wen_60 ? _GEN_7936 : data_0_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7969 = wen_60 ? _GEN_7937 : data_1_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7970 = wen_60 ? _GEN_7938 : data_2_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7971 = wen_60 ? _GEN_7939 : data_3_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7972 = wen_60 ? _GEN_7940 : data_4_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7973 = wen_60 ? _GEN_7941 : data_5_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7974 = wen_60 ? _GEN_7942 : data_6_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7975 = wen_60 ? _GEN_7943 : data_7_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7976 = wen_60 ? _GEN_7944 : data_8_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7977 = wen_60 ? _GEN_7945 : data_9_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7978 = wen_60 ? _GEN_7946 : data_10_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7979 = wen_60 ? _GEN_7947 : data_11_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7980 = wen_60 ? _GEN_7948 : data_12_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7981 = wen_60 ? _GEN_7949 : data_13_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7982 = wen_60 ? _GEN_7950 : data_14_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_7983 = wen_60 ? _GEN_7951 : data_15_7_4; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_7984 = wen_60 ? _GEN_7952 : _GEN_4032; // @[Sbuffer.scala 160:18]
  wire  _GEN_7985 = wen_60 ? _GEN_7953 : _GEN_4033; // @[Sbuffer.scala 160:18]
  wire  _GEN_7986 = wen_60 ? _GEN_7954 : _GEN_4034; // @[Sbuffer.scala 160:18]
  wire  _GEN_7987 = wen_60 ? _GEN_7955 : _GEN_4035; // @[Sbuffer.scala 160:18]
  wire  _GEN_7988 = wen_60 ? _GEN_7956 : _GEN_4036; // @[Sbuffer.scala 160:18]
  wire  _GEN_7989 = wen_60 ? _GEN_7957 : _GEN_4037; // @[Sbuffer.scala 160:18]
  wire  _GEN_7990 = wen_60 ? _GEN_7958 : _GEN_4038; // @[Sbuffer.scala 160:18]
  wire  _GEN_7991 = wen_60 ? _GEN_7959 : _GEN_4039; // @[Sbuffer.scala 160:18]
  wire  _GEN_7992 = wen_60 ? _GEN_7960 : _GEN_4040; // @[Sbuffer.scala 160:18]
  wire  _GEN_7993 = wen_60 ? _GEN_7961 : _GEN_4041; // @[Sbuffer.scala 160:18]
  wire  _GEN_7994 = wen_60 ? _GEN_7962 : _GEN_4042; // @[Sbuffer.scala 160:18]
  wire  _GEN_7995 = wen_60 ? _GEN_7963 : _GEN_4043; // @[Sbuffer.scala 160:18]
  wire  _GEN_7996 = wen_60 ? _GEN_7964 : _GEN_4044; // @[Sbuffer.scala 160:18]
  wire  _GEN_7997 = wen_60 ? _GEN_7965 : _GEN_4045; // @[Sbuffer.scala 160:18]
  wire  _GEN_7998 = wen_60 ? _GEN_7966 : _GEN_4046; // @[Sbuffer.scala 160:18]
  wire  _GEN_7999 = wen_60 ? _GEN_7967 : _GEN_4047; // @[Sbuffer.scala 160:18]
  wire  _wen_T_247 = w_mask_s1_0[5] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_61 = w_valid_s1_0 & _wen_T_247; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_8000 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_0_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8001 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_1_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8002 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_2_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8003 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_3_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8004 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_4_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8005 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_5_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8006 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_6_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8007 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_7_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8008 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_8_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8009 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[47:40] : data_9_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8010 = 4'ha == w_addr_s1_0 ? w_data_s1_0[47:40] : data_10_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8011 = 4'hb == w_addr_s1_0 ? w_data_s1_0[47:40] : data_11_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8012 = 4'hc == w_addr_s1_0 ? w_data_s1_0[47:40] : data_12_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8013 = 4'hd == w_addr_s1_0 ? w_data_s1_0[47:40] : data_13_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8014 = 4'he == w_addr_s1_0 ? w_data_s1_0[47:40] : data_14_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8015 = 4'hf == w_addr_s1_0 ? w_data_s1_0[47:40] : data_15_7_5; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_8016 = 4'h0 == w_addr_s1_0 | _GEN_4048; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8017 = 4'h1 == w_addr_s1_0 | _GEN_4049; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8018 = 4'h2 == w_addr_s1_0 | _GEN_4050; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8019 = 4'h3 == w_addr_s1_0 | _GEN_4051; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8020 = 4'h4 == w_addr_s1_0 | _GEN_4052; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8021 = 4'h5 == w_addr_s1_0 | _GEN_4053; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8022 = 4'h6 == w_addr_s1_0 | _GEN_4054; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8023 = 4'h7 == w_addr_s1_0 | _GEN_4055; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8024 = 4'h8 == w_addr_s1_0 | _GEN_4056; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8025 = 4'h9 == w_addr_s1_0 | _GEN_4057; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8026 = 4'ha == w_addr_s1_0 | _GEN_4058; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8027 = 4'hb == w_addr_s1_0 | _GEN_4059; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8028 = 4'hc == w_addr_s1_0 | _GEN_4060; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8029 = 4'hd == w_addr_s1_0 | _GEN_4061; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8030 = 4'he == w_addr_s1_0 | _GEN_4062; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8031 = 4'hf == w_addr_s1_0 | _GEN_4063; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_8032 = wen_61 ? _GEN_8000 : data_0_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8033 = wen_61 ? _GEN_8001 : data_1_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8034 = wen_61 ? _GEN_8002 : data_2_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8035 = wen_61 ? _GEN_8003 : data_3_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8036 = wen_61 ? _GEN_8004 : data_4_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8037 = wen_61 ? _GEN_8005 : data_5_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8038 = wen_61 ? _GEN_8006 : data_6_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8039 = wen_61 ? _GEN_8007 : data_7_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8040 = wen_61 ? _GEN_8008 : data_8_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8041 = wen_61 ? _GEN_8009 : data_9_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8042 = wen_61 ? _GEN_8010 : data_10_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8043 = wen_61 ? _GEN_8011 : data_11_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8044 = wen_61 ? _GEN_8012 : data_12_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8045 = wen_61 ? _GEN_8013 : data_13_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8046 = wen_61 ? _GEN_8014 : data_14_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8047 = wen_61 ? _GEN_8015 : data_15_7_5; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_8048 = wen_61 ? _GEN_8016 : _GEN_4048; // @[Sbuffer.scala 160:18]
  wire  _GEN_8049 = wen_61 ? _GEN_8017 : _GEN_4049; // @[Sbuffer.scala 160:18]
  wire  _GEN_8050 = wen_61 ? _GEN_8018 : _GEN_4050; // @[Sbuffer.scala 160:18]
  wire  _GEN_8051 = wen_61 ? _GEN_8019 : _GEN_4051; // @[Sbuffer.scala 160:18]
  wire  _GEN_8052 = wen_61 ? _GEN_8020 : _GEN_4052; // @[Sbuffer.scala 160:18]
  wire  _GEN_8053 = wen_61 ? _GEN_8021 : _GEN_4053; // @[Sbuffer.scala 160:18]
  wire  _GEN_8054 = wen_61 ? _GEN_8022 : _GEN_4054; // @[Sbuffer.scala 160:18]
  wire  _GEN_8055 = wen_61 ? _GEN_8023 : _GEN_4055; // @[Sbuffer.scala 160:18]
  wire  _GEN_8056 = wen_61 ? _GEN_8024 : _GEN_4056; // @[Sbuffer.scala 160:18]
  wire  _GEN_8057 = wen_61 ? _GEN_8025 : _GEN_4057; // @[Sbuffer.scala 160:18]
  wire  _GEN_8058 = wen_61 ? _GEN_8026 : _GEN_4058; // @[Sbuffer.scala 160:18]
  wire  _GEN_8059 = wen_61 ? _GEN_8027 : _GEN_4059; // @[Sbuffer.scala 160:18]
  wire  _GEN_8060 = wen_61 ? _GEN_8028 : _GEN_4060; // @[Sbuffer.scala 160:18]
  wire  _GEN_8061 = wen_61 ? _GEN_8029 : _GEN_4061; // @[Sbuffer.scala 160:18]
  wire  _GEN_8062 = wen_61 ? _GEN_8030 : _GEN_4062; // @[Sbuffer.scala 160:18]
  wire  _GEN_8063 = wen_61 ? _GEN_8031 : _GEN_4063; // @[Sbuffer.scala 160:18]
  wire  _wen_T_251 = w_mask_s1_0[6] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_62 = w_valid_s1_0 & _wen_T_251; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_8064 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_0_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8065 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_1_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8066 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_2_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8067 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_3_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8068 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_4_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8069 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_5_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8070 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_6_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8071 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_7_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8072 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_8_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8073 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[55:48] : data_9_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8074 = 4'ha == w_addr_s1_0 ? w_data_s1_0[55:48] : data_10_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8075 = 4'hb == w_addr_s1_0 ? w_data_s1_0[55:48] : data_11_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8076 = 4'hc == w_addr_s1_0 ? w_data_s1_0[55:48] : data_12_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8077 = 4'hd == w_addr_s1_0 ? w_data_s1_0[55:48] : data_13_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8078 = 4'he == w_addr_s1_0 ? w_data_s1_0[55:48] : data_14_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8079 = 4'hf == w_addr_s1_0 ? w_data_s1_0[55:48] : data_15_7_6; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_8080 = 4'h0 == w_addr_s1_0 | _GEN_4064; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8081 = 4'h1 == w_addr_s1_0 | _GEN_4065; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8082 = 4'h2 == w_addr_s1_0 | _GEN_4066; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8083 = 4'h3 == w_addr_s1_0 | _GEN_4067; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8084 = 4'h4 == w_addr_s1_0 | _GEN_4068; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8085 = 4'h5 == w_addr_s1_0 | _GEN_4069; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8086 = 4'h6 == w_addr_s1_0 | _GEN_4070; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8087 = 4'h7 == w_addr_s1_0 | _GEN_4071; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8088 = 4'h8 == w_addr_s1_0 | _GEN_4072; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8089 = 4'h9 == w_addr_s1_0 | _GEN_4073; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8090 = 4'ha == w_addr_s1_0 | _GEN_4074; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8091 = 4'hb == w_addr_s1_0 | _GEN_4075; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8092 = 4'hc == w_addr_s1_0 | _GEN_4076; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8093 = 4'hd == w_addr_s1_0 | _GEN_4077; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8094 = 4'he == w_addr_s1_0 | _GEN_4078; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8095 = 4'hf == w_addr_s1_0 | _GEN_4079; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_8096 = wen_62 ? _GEN_8064 : data_0_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8097 = wen_62 ? _GEN_8065 : data_1_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8098 = wen_62 ? _GEN_8066 : data_2_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8099 = wen_62 ? _GEN_8067 : data_3_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8100 = wen_62 ? _GEN_8068 : data_4_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8101 = wen_62 ? _GEN_8069 : data_5_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8102 = wen_62 ? _GEN_8070 : data_6_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8103 = wen_62 ? _GEN_8071 : data_7_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8104 = wen_62 ? _GEN_8072 : data_8_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8105 = wen_62 ? _GEN_8073 : data_9_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8106 = wen_62 ? _GEN_8074 : data_10_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8107 = wen_62 ? _GEN_8075 : data_11_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8108 = wen_62 ? _GEN_8076 : data_12_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8109 = wen_62 ? _GEN_8077 : data_13_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8110 = wen_62 ? _GEN_8078 : data_14_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8111 = wen_62 ? _GEN_8079 : data_15_7_6; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_8112 = wen_62 ? _GEN_8080 : _GEN_4064; // @[Sbuffer.scala 160:18]
  wire  _GEN_8113 = wen_62 ? _GEN_8081 : _GEN_4065; // @[Sbuffer.scala 160:18]
  wire  _GEN_8114 = wen_62 ? _GEN_8082 : _GEN_4066; // @[Sbuffer.scala 160:18]
  wire  _GEN_8115 = wen_62 ? _GEN_8083 : _GEN_4067; // @[Sbuffer.scala 160:18]
  wire  _GEN_8116 = wen_62 ? _GEN_8084 : _GEN_4068; // @[Sbuffer.scala 160:18]
  wire  _GEN_8117 = wen_62 ? _GEN_8085 : _GEN_4069; // @[Sbuffer.scala 160:18]
  wire  _GEN_8118 = wen_62 ? _GEN_8086 : _GEN_4070; // @[Sbuffer.scala 160:18]
  wire  _GEN_8119 = wen_62 ? _GEN_8087 : _GEN_4071; // @[Sbuffer.scala 160:18]
  wire  _GEN_8120 = wen_62 ? _GEN_8088 : _GEN_4072; // @[Sbuffer.scala 160:18]
  wire  _GEN_8121 = wen_62 ? _GEN_8089 : _GEN_4073; // @[Sbuffer.scala 160:18]
  wire  _GEN_8122 = wen_62 ? _GEN_8090 : _GEN_4074; // @[Sbuffer.scala 160:18]
  wire  _GEN_8123 = wen_62 ? _GEN_8091 : _GEN_4075; // @[Sbuffer.scala 160:18]
  wire  _GEN_8124 = wen_62 ? _GEN_8092 : _GEN_4076; // @[Sbuffer.scala 160:18]
  wire  _GEN_8125 = wen_62 ? _GEN_8093 : _GEN_4077; // @[Sbuffer.scala 160:18]
  wire  _GEN_8126 = wen_62 ? _GEN_8094 : _GEN_4078; // @[Sbuffer.scala 160:18]
  wire  _GEN_8127 = wen_62 ? _GEN_8095 : _GEN_4079; // @[Sbuffer.scala 160:18]
  wire  _wen_T_255 = w_mask_s1_0[7] & w_word_offset_s1_0 == 3'h7 | w_wline_s1_0; // @[Sbuffer.scala 157:70]
  wire  wen_63 = w_valid_s1_0 & _wen_T_255; // @[Sbuffer.scala 156:25]
  wire [7:0] _GEN_8128 = 4'h0 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_0_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8129 = 4'h1 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_1_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8130 = 4'h2 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_2_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8131 = 4'h3 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_3_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8132 = 4'h4 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_4_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8133 = 4'h5 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_5_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8134 = 4'h6 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_6_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8135 = 4'h7 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_7_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8136 = 4'h8 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_8_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8137 = 4'h9 == w_addr_s1_0 ? w_data_s1_0[63:56] : data_9_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8138 = 4'ha == w_addr_s1_0 ? w_data_s1_0[63:56] : data_10_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8139 = 4'hb == w_addr_s1_0 ? w_data_s1_0[63:56] : data_11_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8140 = 4'hc == w_addr_s1_0 ? w_data_s1_0[63:56] : data_12_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8141 = 4'hd == w_addr_s1_0 ? w_data_s1_0[63:56] : data_13_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8142 = 4'he == w_addr_s1_0 ? w_data_s1_0[63:56] : data_14_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire [7:0] _GEN_8143 = 4'hf == w_addr_s1_0 ? w_data_s1_0[63:56] : data_15_7_7; // @[Sbuffer.scala 161:{42,42} 96:17]
  wire  _GEN_8144 = 4'h0 == w_addr_s1_0 | _GEN_4080; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8145 = 4'h1 == w_addr_s1_0 | _GEN_4081; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8146 = 4'h2 == w_addr_s1_0 | _GEN_4082; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8147 = 4'h3 == w_addr_s1_0 | _GEN_4083; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8148 = 4'h4 == w_addr_s1_0 | _GEN_4084; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8149 = 4'h5 == w_addr_s1_0 | _GEN_4085; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8150 = 4'h6 == w_addr_s1_0 | _GEN_4086; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8151 = 4'h7 == w_addr_s1_0 | _GEN_4087; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8152 = 4'h8 == w_addr_s1_0 | _GEN_4088; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8153 = 4'h9 == w_addr_s1_0 | _GEN_4089; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8154 = 4'ha == w_addr_s1_0 | _GEN_4090; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8155 = 4'hb == w_addr_s1_0 | _GEN_4091; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8156 = 4'hc == w_addr_s1_0 | _GEN_4092; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8157 = 4'hd == w_addr_s1_0 | _GEN_4093; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8158 = 4'he == w_addr_s1_0 | _GEN_4094; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8159 = 4'hf == w_addr_s1_0 | _GEN_4095; // @[Sbuffer.scala 162:{42,42}]
  wire [7:0] _GEN_8160 = wen_63 ? _GEN_8128 : data_0_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8161 = wen_63 ? _GEN_8129 : data_1_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8162 = wen_63 ? _GEN_8130 : data_2_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8163 = wen_63 ? _GEN_8131 : data_3_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8164 = wen_63 ? _GEN_8132 : data_4_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8165 = wen_63 ? _GEN_8133 : data_5_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8166 = wen_63 ? _GEN_8134 : data_6_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8167 = wen_63 ? _GEN_8135 : data_7_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8168 = wen_63 ? _GEN_8136 : data_8_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8169 = wen_63 ? _GEN_8137 : data_9_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8170 = wen_63 ? _GEN_8138 : data_10_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8171 = wen_63 ? _GEN_8139 : data_11_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8172 = wen_63 ? _GEN_8140 : data_12_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8173 = wen_63 ? _GEN_8141 : data_13_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8174 = wen_63 ? _GEN_8142 : data_14_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire [7:0] _GEN_8175 = wen_63 ? _GEN_8143 : data_15_7_7; // @[Sbuffer.scala 160:18 96:17]
  wire  _GEN_8176 = wen_63 ? _GEN_8144 : _GEN_4080; // @[Sbuffer.scala 160:18]
  wire  _GEN_8177 = wen_63 ? _GEN_8145 : _GEN_4081; // @[Sbuffer.scala 160:18]
  wire  _GEN_8178 = wen_63 ? _GEN_8146 : _GEN_4082; // @[Sbuffer.scala 160:18]
  wire  _GEN_8179 = wen_63 ? _GEN_8147 : _GEN_4083; // @[Sbuffer.scala 160:18]
  wire  _GEN_8180 = wen_63 ? _GEN_8148 : _GEN_4084; // @[Sbuffer.scala 160:18]
  wire  _GEN_8181 = wen_63 ? _GEN_8149 : _GEN_4085; // @[Sbuffer.scala 160:18]
  wire  _GEN_8182 = wen_63 ? _GEN_8150 : _GEN_4086; // @[Sbuffer.scala 160:18]
  wire  _GEN_8183 = wen_63 ? _GEN_8151 : _GEN_4087; // @[Sbuffer.scala 160:18]
  wire  _GEN_8184 = wen_63 ? _GEN_8152 : _GEN_4088; // @[Sbuffer.scala 160:18]
  wire  _GEN_8185 = wen_63 ? _GEN_8153 : _GEN_4089; // @[Sbuffer.scala 160:18]
  wire  _GEN_8186 = wen_63 ? _GEN_8154 : _GEN_4090; // @[Sbuffer.scala 160:18]
  wire  _GEN_8187 = wen_63 ? _GEN_8155 : _GEN_4091; // @[Sbuffer.scala 160:18]
  wire  _GEN_8188 = wen_63 ? _GEN_8156 : _GEN_4092; // @[Sbuffer.scala 160:18]
  wire  _GEN_8189 = wen_63 ? _GEN_8157 : _GEN_4093; // @[Sbuffer.scala 160:18]
  wire  _GEN_8190 = wen_63 ? _GEN_8158 : _GEN_4094; // @[Sbuffer.scala 160:18]
  wire  _GEN_8191 = wen_63 ? _GEN_8159 : _GEN_4095; // @[Sbuffer.scala 160:18]
  wire  _wen_T_259 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_64 = w_valid_s1_1 & _wen_T_259; // @[Sbuffer.scala 156:25]
  wire  _GEN_8208 = 4'h0 == w_addr_s1_1 | _GEN_4144; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8209 = 4'h1 == w_addr_s1_1 | _GEN_4145; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8210 = 4'h2 == w_addr_s1_1 | _GEN_4146; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8211 = 4'h3 == w_addr_s1_1 | _GEN_4147; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8212 = 4'h4 == w_addr_s1_1 | _GEN_4148; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8213 = 4'h5 == w_addr_s1_1 | _GEN_4149; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8214 = 4'h6 == w_addr_s1_1 | _GEN_4150; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8215 = 4'h7 == w_addr_s1_1 | _GEN_4151; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8216 = 4'h8 == w_addr_s1_1 | _GEN_4152; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8217 = 4'h9 == w_addr_s1_1 | _GEN_4153; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8218 = 4'ha == w_addr_s1_1 | _GEN_4154; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8219 = 4'hb == w_addr_s1_1 | _GEN_4155; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8220 = 4'hc == w_addr_s1_1 | _GEN_4156; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8221 = 4'hd == w_addr_s1_1 | _GEN_4157; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8222 = 4'he == w_addr_s1_1 | _GEN_4158; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8223 = 4'hf == w_addr_s1_1 | _GEN_4159; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_263 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_65 = w_valid_s1_1 & _wen_T_263; // @[Sbuffer.scala 156:25]
  wire  _GEN_8272 = 4'h0 == w_addr_s1_1 | _GEN_4208; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8273 = 4'h1 == w_addr_s1_1 | _GEN_4209; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8274 = 4'h2 == w_addr_s1_1 | _GEN_4210; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8275 = 4'h3 == w_addr_s1_1 | _GEN_4211; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8276 = 4'h4 == w_addr_s1_1 | _GEN_4212; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8277 = 4'h5 == w_addr_s1_1 | _GEN_4213; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8278 = 4'h6 == w_addr_s1_1 | _GEN_4214; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8279 = 4'h7 == w_addr_s1_1 | _GEN_4215; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8280 = 4'h8 == w_addr_s1_1 | _GEN_4216; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8281 = 4'h9 == w_addr_s1_1 | _GEN_4217; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8282 = 4'ha == w_addr_s1_1 | _GEN_4218; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8283 = 4'hb == w_addr_s1_1 | _GEN_4219; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8284 = 4'hc == w_addr_s1_1 | _GEN_4220; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8285 = 4'hd == w_addr_s1_1 | _GEN_4221; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8286 = 4'he == w_addr_s1_1 | _GEN_4222; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8287 = 4'hf == w_addr_s1_1 | _GEN_4223; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_267 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_66 = w_valid_s1_1 & _wen_T_267; // @[Sbuffer.scala 156:25]
  wire  _GEN_8336 = 4'h0 == w_addr_s1_1 | _GEN_4272; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8337 = 4'h1 == w_addr_s1_1 | _GEN_4273; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8338 = 4'h2 == w_addr_s1_1 | _GEN_4274; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8339 = 4'h3 == w_addr_s1_1 | _GEN_4275; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8340 = 4'h4 == w_addr_s1_1 | _GEN_4276; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8341 = 4'h5 == w_addr_s1_1 | _GEN_4277; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8342 = 4'h6 == w_addr_s1_1 | _GEN_4278; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8343 = 4'h7 == w_addr_s1_1 | _GEN_4279; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8344 = 4'h8 == w_addr_s1_1 | _GEN_4280; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8345 = 4'h9 == w_addr_s1_1 | _GEN_4281; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8346 = 4'ha == w_addr_s1_1 | _GEN_4282; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8347 = 4'hb == w_addr_s1_1 | _GEN_4283; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8348 = 4'hc == w_addr_s1_1 | _GEN_4284; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8349 = 4'hd == w_addr_s1_1 | _GEN_4285; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8350 = 4'he == w_addr_s1_1 | _GEN_4286; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8351 = 4'hf == w_addr_s1_1 | _GEN_4287; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_271 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_67 = w_valid_s1_1 & _wen_T_271; // @[Sbuffer.scala 156:25]
  wire  _GEN_8400 = 4'h0 == w_addr_s1_1 | _GEN_4336; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8401 = 4'h1 == w_addr_s1_1 | _GEN_4337; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8402 = 4'h2 == w_addr_s1_1 | _GEN_4338; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8403 = 4'h3 == w_addr_s1_1 | _GEN_4339; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8404 = 4'h4 == w_addr_s1_1 | _GEN_4340; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8405 = 4'h5 == w_addr_s1_1 | _GEN_4341; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8406 = 4'h6 == w_addr_s1_1 | _GEN_4342; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8407 = 4'h7 == w_addr_s1_1 | _GEN_4343; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8408 = 4'h8 == w_addr_s1_1 | _GEN_4344; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8409 = 4'h9 == w_addr_s1_1 | _GEN_4345; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8410 = 4'ha == w_addr_s1_1 | _GEN_4346; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8411 = 4'hb == w_addr_s1_1 | _GEN_4347; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8412 = 4'hc == w_addr_s1_1 | _GEN_4348; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8413 = 4'hd == w_addr_s1_1 | _GEN_4349; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8414 = 4'he == w_addr_s1_1 | _GEN_4350; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8415 = 4'hf == w_addr_s1_1 | _GEN_4351; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_275 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_68 = w_valid_s1_1 & _wen_T_275; // @[Sbuffer.scala 156:25]
  wire  _GEN_8464 = 4'h0 == w_addr_s1_1 | _GEN_4400; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8465 = 4'h1 == w_addr_s1_1 | _GEN_4401; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8466 = 4'h2 == w_addr_s1_1 | _GEN_4402; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8467 = 4'h3 == w_addr_s1_1 | _GEN_4403; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8468 = 4'h4 == w_addr_s1_1 | _GEN_4404; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8469 = 4'h5 == w_addr_s1_1 | _GEN_4405; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8470 = 4'h6 == w_addr_s1_1 | _GEN_4406; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8471 = 4'h7 == w_addr_s1_1 | _GEN_4407; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8472 = 4'h8 == w_addr_s1_1 | _GEN_4408; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8473 = 4'h9 == w_addr_s1_1 | _GEN_4409; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8474 = 4'ha == w_addr_s1_1 | _GEN_4410; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8475 = 4'hb == w_addr_s1_1 | _GEN_4411; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8476 = 4'hc == w_addr_s1_1 | _GEN_4412; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8477 = 4'hd == w_addr_s1_1 | _GEN_4413; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8478 = 4'he == w_addr_s1_1 | _GEN_4414; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8479 = 4'hf == w_addr_s1_1 | _GEN_4415; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_279 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_69 = w_valid_s1_1 & _wen_T_279; // @[Sbuffer.scala 156:25]
  wire  _GEN_8528 = 4'h0 == w_addr_s1_1 | _GEN_4464; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8529 = 4'h1 == w_addr_s1_1 | _GEN_4465; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8530 = 4'h2 == w_addr_s1_1 | _GEN_4466; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8531 = 4'h3 == w_addr_s1_1 | _GEN_4467; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8532 = 4'h4 == w_addr_s1_1 | _GEN_4468; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8533 = 4'h5 == w_addr_s1_1 | _GEN_4469; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8534 = 4'h6 == w_addr_s1_1 | _GEN_4470; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8535 = 4'h7 == w_addr_s1_1 | _GEN_4471; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8536 = 4'h8 == w_addr_s1_1 | _GEN_4472; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8537 = 4'h9 == w_addr_s1_1 | _GEN_4473; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8538 = 4'ha == w_addr_s1_1 | _GEN_4474; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8539 = 4'hb == w_addr_s1_1 | _GEN_4475; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8540 = 4'hc == w_addr_s1_1 | _GEN_4476; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8541 = 4'hd == w_addr_s1_1 | _GEN_4477; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8542 = 4'he == w_addr_s1_1 | _GEN_4478; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8543 = 4'hf == w_addr_s1_1 | _GEN_4479; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_283 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_70 = w_valid_s1_1 & _wen_T_283; // @[Sbuffer.scala 156:25]
  wire  _GEN_8592 = 4'h0 == w_addr_s1_1 | _GEN_4528; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8593 = 4'h1 == w_addr_s1_1 | _GEN_4529; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8594 = 4'h2 == w_addr_s1_1 | _GEN_4530; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8595 = 4'h3 == w_addr_s1_1 | _GEN_4531; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8596 = 4'h4 == w_addr_s1_1 | _GEN_4532; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8597 = 4'h5 == w_addr_s1_1 | _GEN_4533; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8598 = 4'h6 == w_addr_s1_1 | _GEN_4534; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8599 = 4'h7 == w_addr_s1_1 | _GEN_4535; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8600 = 4'h8 == w_addr_s1_1 | _GEN_4536; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8601 = 4'h9 == w_addr_s1_1 | _GEN_4537; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8602 = 4'ha == w_addr_s1_1 | _GEN_4538; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8603 = 4'hb == w_addr_s1_1 | _GEN_4539; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8604 = 4'hc == w_addr_s1_1 | _GEN_4540; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8605 = 4'hd == w_addr_s1_1 | _GEN_4541; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8606 = 4'he == w_addr_s1_1 | _GEN_4542; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8607 = 4'hf == w_addr_s1_1 | _GEN_4543; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_287 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h0 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_71 = w_valid_s1_1 & _wen_T_287; // @[Sbuffer.scala 156:25]
  wire  _GEN_8656 = 4'h0 == w_addr_s1_1 | _GEN_4592; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8657 = 4'h1 == w_addr_s1_1 | _GEN_4593; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8658 = 4'h2 == w_addr_s1_1 | _GEN_4594; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8659 = 4'h3 == w_addr_s1_1 | _GEN_4595; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8660 = 4'h4 == w_addr_s1_1 | _GEN_4596; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8661 = 4'h5 == w_addr_s1_1 | _GEN_4597; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8662 = 4'h6 == w_addr_s1_1 | _GEN_4598; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8663 = 4'h7 == w_addr_s1_1 | _GEN_4599; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8664 = 4'h8 == w_addr_s1_1 | _GEN_4600; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8665 = 4'h9 == w_addr_s1_1 | _GEN_4601; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8666 = 4'ha == w_addr_s1_1 | _GEN_4602; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8667 = 4'hb == w_addr_s1_1 | _GEN_4603; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8668 = 4'hc == w_addr_s1_1 | _GEN_4604; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8669 = 4'hd == w_addr_s1_1 | _GEN_4605; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8670 = 4'he == w_addr_s1_1 | _GEN_4606; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8671 = 4'hf == w_addr_s1_1 | _GEN_4607; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_291 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_72 = w_valid_s1_1 & _wen_T_291; // @[Sbuffer.scala 156:25]
  wire  _GEN_8720 = 4'h0 == w_addr_s1_1 | _GEN_4656; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8721 = 4'h1 == w_addr_s1_1 | _GEN_4657; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8722 = 4'h2 == w_addr_s1_1 | _GEN_4658; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8723 = 4'h3 == w_addr_s1_1 | _GEN_4659; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8724 = 4'h4 == w_addr_s1_1 | _GEN_4660; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8725 = 4'h5 == w_addr_s1_1 | _GEN_4661; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8726 = 4'h6 == w_addr_s1_1 | _GEN_4662; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8727 = 4'h7 == w_addr_s1_1 | _GEN_4663; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8728 = 4'h8 == w_addr_s1_1 | _GEN_4664; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8729 = 4'h9 == w_addr_s1_1 | _GEN_4665; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8730 = 4'ha == w_addr_s1_1 | _GEN_4666; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8731 = 4'hb == w_addr_s1_1 | _GEN_4667; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8732 = 4'hc == w_addr_s1_1 | _GEN_4668; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8733 = 4'hd == w_addr_s1_1 | _GEN_4669; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8734 = 4'he == w_addr_s1_1 | _GEN_4670; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8735 = 4'hf == w_addr_s1_1 | _GEN_4671; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_295 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_73 = w_valid_s1_1 & _wen_T_295; // @[Sbuffer.scala 156:25]
  wire  _GEN_8784 = 4'h0 == w_addr_s1_1 | _GEN_4720; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8785 = 4'h1 == w_addr_s1_1 | _GEN_4721; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8786 = 4'h2 == w_addr_s1_1 | _GEN_4722; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8787 = 4'h3 == w_addr_s1_1 | _GEN_4723; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8788 = 4'h4 == w_addr_s1_1 | _GEN_4724; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8789 = 4'h5 == w_addr_s1_1 | _GEN_4725; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8790 = 4'h6 == w_addr_s1_1 | _GEN_4726; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8791 = 4'h7 == w_addr_s1_1 | _GEN_4727; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8792 = 4'h8 == w_addr_s1_1 | _GEN_4728; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8793 = 4'h9 == w_addr_s1_1 | _GEN_4729; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8794 = 4'ha == w_addr_s1_1 | _GEN_4730; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8795 = 4'hb == w_addr_s1_1 | _GEN_4731; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8796 = 4'hc == w_addr_s1_1 | _GEN_4732; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8797 = 4'hd == w_addr_s1_1 | _GEN_4733; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8798 = 4'he == w_addr_s1_1 | _GEN_4734; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8799 = 4'hf == w_addr_s1_1 | _GEN_4735; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_299 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_74 = w_valid_s1_1 & _wen_T_299; // @[Sbuffer.scala 156:25]
  wire  _GEN_8848 = 4'h0 == w_addr_s1_1 | _GEN_4784; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8849 = 4'h1 == w_addr_s1_1 | _GEN_4785; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8850 = 4'h2 == w_addr_s1_1 | _GEN_4786; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8851 = 4'h3 == w_addr_s1_1 | _GEN_4787; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8852 = 4'h4 == w_addr_s1_1 | _GEN_4788; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8853 = 4'h5 == w_addr_s1_1 | _GEN_4789; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8854 = 4'h6 == w_addr_s1_1 | _GEN_4790; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8855 = 4'h7 == w_addr_s1_1 | _GEN_4791; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8856 = 4'h8 == w_addr_s1_1 | _GEN_4792; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8857 = 4'h9 == w_addr_s1_1 | _GEN_4793; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8858 = 4'ha == w_addr_s1_1 | _GEN_4794; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8859 = 4'hb == w_addr_s1_1 | _GEN_4795; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8860 = 4'hc == w_addr_s1_1 | _GEN_4796; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8861 = 4'hd == w_addr_s1_1 | _GEN_4797; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8862 = 4'he == w_addr_s1_1 | _GEN_4798; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8863 = 4'hf == w_addr_s1_1 | _GEN_4799; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_303 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_75 = w_valid_s1_1 & _wen_T_303; // @[Sbuffer.scala 156:25]
  wire  _GEN_8912 = 4'h0 == w_addr_s1_1 | _GEN_4848; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8913 = 4'h1 == w_addr_s1_1 | _GEN_4849; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8914 = 4'h2 == w_addr_s1_1 | _GEN_4850; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8915 = 4'h3 == w_addr_s1_1 | _GEN_4851; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8916 = 4'h4 == w_addr_s1_1 | _GEN_4852; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8917 = 4'h5 == w_addr_s1_1 | _GEN_4853; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8918 = 4'h6 == w_addr_s1_1 | _GEN_4854; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8919 = 4'h7 == w_addr_s1_1 | _GEN_4855; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8920 = 4'h8 == w_addr_s1_1 | _GEN_4856; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8921 = 4'h9 == w_addr_s1_1 | _GEN_4857; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8922 = 4'ha == w_addr_s1_1 | _GEN_4858; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8923 = 4'hb == w_addr_s1_1 | _GEN_4859; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8924 = 4'hc == w_addr_s1_1 | _GEN_4860; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8925 = 4'hd == w_addr_s1_1 | _GEN_4861; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8926 = 4'he == w_addr_s1_1 | _GEN_4862; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8927 = 4'hf == w_addr_s1_1 | _GEN_4863; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_307 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_76 = w_valid_s1_1 & _wen_T_307; // @[Sbuffer.scala 156:25]
  wire  _GEN_8976 = 4'h0 == w_addr_s1_1 | _GEN_4912; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8977 = 4'h1 == w_addr_s1_1 | _GEN_4913; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8978 = 4'h2 == w_addr_s1_1 | _GEN_4914; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8979 = 4'h3 == w_addr_s1_1 | _GEN_4915; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8980 = 4'h4 == w_addr_s1_1 | _GEN_4916; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8981 = 4'h5 == w_addr_s1_1 | _GEN_4917; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8982 = 4'h6 == w_addr_s1_1 | _GEN_4918; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8983 = 4'h7 == w_addr_s1_1 | _GEN_4919; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8984 = 4'h8 == w_addr_s1_1 | _GEN_4920; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8985 = 4'h9 == w_addr_s1_1 | _GEN_4921; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8986 = 4'ha == w_addr_s1_1 | _GEN_4922; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8987 = 4'hb == w_addr_s1_1 | _GEN_4923; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8988 = 4'hc == w_addr_s1_1 | _GEN_4924; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8989 = 4'hd == w_addr_s1_1 | _GEN_4925; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8990 = 4'he == w_addr_s1_1 | _GEN_4926; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_8991 = 4'hf == w_addr_s1_1 | _GEN_4927; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_311 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_77 = w_valid_s1_1 & _wen_T_311; // @[Sbuffer.scala 156:25]
  wire  _GEN_9040 = 4'h0 == w_addr_s1_1 | _GEN_4976; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9041 = 4'h1 == w_addr_s1_1 | _GEN_4977; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9042 = 4'h2 == w_addr_s1_1 | _GEN_4978; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9043 = 4'h3 == w_addr_s1_1 | _GEN_4979; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9044 = 4'h4 == w_addr_s1_1 | _GEN_4980; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9045 = 4'h5 == w_addr_s1_1 | _GEN_4981; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9046 = 4'h6 == w_addr_s1_1 | _GEN_4982; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9047 = 4'h7 == w_addr_s1_1 | _GEN_4983; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9048 = 4'h8 == w_addr_s1_1 | _GEN_4984; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9049 = 4'h9 == w_addr_s1_1 | _GEN_4985; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9050 = 4'ha == w_addr_s1_1 | _GEN_4986; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9051 = 4'hb == w_addr_s1_1 | _GEN_4987; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9052 = 4'hc == w_addr_s1_1 | _GEN_4988; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9053 = 4'hd == w_addr_s1_1 | _GEN_4989; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9054 = 4'he == w_addr_s1_1 | _GEN_4990; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9055 = 4'hf == w_addr_s1_1 | _GEN_4991; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_315 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_78 = w_valid_s1_1 & _wen_T_315; // @[Sbuffer.scala 156:25]
  wire  _GEN_9104 = 4'h0 == w_addr_s1_1 | _GEN_5040; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9105 = 4'h1 == w_addr_s1_1 | _GEN_5041; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9106 = 4'h2 == w_addr_s1_1 | _GEN_5042; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9107 = 4'h3 == w_addr_s1_1 | _GEN_5043; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9108 = 4'h4 == w_addr_s1_1 | _GEN_5044; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9109 = 4'h5 == w_addr_s1_1 | _GEN_5045; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9110 = 4'h6 == w_addr_s1_1 | _GEN_5046; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9111 = 4'h7 == w_addr_s1_1 | _GEN_5047; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9112 = 4'h8 == w_addr_s1_1 | _GEN_5048; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9113 = 4'h9 == w_addr_s1_1 | _GEN_5049; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9114 = 4'ha == w_addr_s1_1 | _GEN_5050; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9115 = 4'hb == w_addr_s1_1 | _GEN_5051; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9116 = 4'hc == w_addr_s1_1 | _GEN_5052; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9117 = 4'hd == w_addr_s1_1 | _GEN_5053; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9118 = 4'he == w_addr_s1_1 | _GEN_5054; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9119 = 4'hf == w_addr_s1_1 | _GEN_5055; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_319 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h1 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_79 = w_valid_s1_1 & _wen_T_319; // @[Sbuffer.scala 156:25]
  wire  _GEN_9168 = 4'h0 == w_addr_s1_1 | _GEN_5104; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9169 = 4'h1 == w_addr_s1_1 | _GEN_5105; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9170 = 4'h2 == w_addr_s1_1 | _GEN_5106; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9171 = 4'h3 == w_addr_s1_1 | _GEN_5107; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9172 = 4'h4 == w_addr_s1_1 | _GEN_5108; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9173 = 4'h5 == w_addr_s1_1 | _GEN_5109; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9174 = 4'h6 == w_addr_s1_1 | _GEN_5110; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9175 = 4'h7 == w_addr_s1_1 | _GEN_5111; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9176 = 4'h8 == w_addr_s1_1 | _GEN_5112; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9177 = 4'h9 == w_addr_s1_1 | _GEN_5113; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9178 = 4'ha == w_addr_s1_1 | _GEN_5114; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9179 = 4'hb == w_addr_s1_1 | _GEN_5115; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9180 = 4'hc == w_addr_s1_1 | _GEN_5116; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9181 = 4'hd == w_addr_s1_1 | _GEN_5117; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9182 = 4'he == w_addr_s1_1 | _GEN_5118; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9183 = 4'hf == w_addr_s1_1 | _GEN_5119; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_323 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_80 = w_valid_s1_1 & _wen_T_323; // @[Sbuffer.scala 156:25]
  wire  _GEN_9232 = 4'h0 == w_addr_s1_1 | _GEN_5168; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9233 = 4'h1 == w_addr_s1_1 | _GEN_5169; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9234 = 4'h2 == w_addr_s1_1 | _GEN_5170; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9235 = 4'h3 == w_addr_s1_1 | _GEN_5171; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9236 = 4'h4 == w_addr_s1_1 | _GEN_5172; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9237 = 4'h5 == w_addr_s1_1 | _GEN_5173; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9238 = 4'h6 == w_addr_s1_1 | _GEN_5174; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9239 = 4'h7 == w_addr_s1_1 | _GEN_5175; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9240 = 4'h8 == w_addr_s1_1 | _GEN_5176; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9241 = 4'h9 == w_addr_s1_1 | _GEN_5177; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9242 = 4'ha == w_addr_s1_1 | _GEN_5178; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9243 = 4'hb == w_addr_s1_1 | _GEN_5179; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9244 = 4'hc == w_addr_s1_1 | _GEN_5180; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9245 = 4'hd == w_addr_s1_1 | _GEN_5181; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9246 = 4'he == w_addr_s1_1 | _GEN_5182; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9247 = 4'hf == w_addr_s1_1 | _GEN_5183; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_327 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_81 = w_valid_s1_1 & _wen_T_327; // @[Sbuffer.scala 156:25]
  wire  _GEN_9296 = 4'h0 == w_addr_s1_1 | _GEN_5232; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9297 = 4'h1 == w_addr_s1_1 | _GEN_5233; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9298 = 4'h2 == w_addr_s1_1 | _GEN_5234; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9299 = 4'h3 == w_addr_s1_1 | _GEN_5235; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9300 = 4'h4 == w_addr_s1_1 | _GEN_5236; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9301 = 4'h5 == w_addr_s1_1 | _GEN_5237; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9302 = 4'h6 == w_addr_s1_1 | _GEN_5238; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9303 = 4'h7 == w_addr_s1_1 | _GEN_5239; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9304 = 4'h8 == w_addr_s1_1 | _GEN_5240; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9305 = 4'h9 == w_addr_s1_1 | _GEN_5241; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9306 = 4'ha == w_addr_s1_1 | _GEN_5242; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9307 = 4'hb == w_addr_s1_1 | _GEN_5243; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9308 = 4'hc == w_addr_s1_1 | _GEN_5244; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9309 = 4'hd == w_addr_s1_1 | _GEN_5245; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9310 = 4'he == w_addr_s1_1 | _GEN_5246; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9311 = 4'hf == w_addr_s1_1 | _GEN_5247; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_331 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_82 = w_valid_s1_1 & _wen_T_331; // @[Sbuffer.scala 156:25]
  wire  _GEN_9360 = 4'h0 == w_addr_s1_1 | _GEN_5296; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9361 = 4'h1 == w_addr_s1_1 | _GEN_5297; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9362 = 4'h2 == w_addr_s1_1 | _GEN_5298; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9363 = 4'h3 == w_addr_s1_1 | _GEN_5299; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9364 = 4'h4 == w_addr_s1_1 | _GEN_5300; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9365 = 4'h5 == w_addr_s1_1 | _GEN_5301; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9366 = 4'h6 == w_addr_s1_1 | _GEN_5302; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9367 = 4'h7 == w_addr_s1_1 | _GEN_5303; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9368 = 4'h8 == w_addr_s1_1 | _GEN_5304; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9369 = 4'h9 == w_addr_s1_1 | _GEN_5305; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9370 = 4'ha == w_addr_s1_1 | _GEN_5306; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9371 = 4'hb == w_addr_s1_1 | _GEN_5307; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9372 = 4'hc == w_addr_s1_1 | _GEN_5308; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9373 = 4'hd == w_addr_s1_1 | _GEN_5309; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9374 = 4'he == w_addr_s1_1 | _GEN_5310; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9375 = 4'hf == w_addr_s1_1 | _GEN_5311; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_335 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_83 = w_valid_s1_1 & _wen_T_335; // @[Sbuffer.scala 156:25]
  wire  _GEN_9424 = 4'h0 == w_addr_s1_1 | _GEN_5360; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9425 = 4'h1 == w_addr_s1_1 | _GEN_5361; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9426 = 4'h2 == w_addr_s1_1 | _GEN_5362; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9427 = 4'h3 == w_addr_s1_1 | _GEN_5363; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9428 = 4'h4 == w_addr_s1_1 | _GEN_5364; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9429 = 4'h5 == w_addr_s1_1 | _GEN_5365; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9430 = 4'h6 == w_addr_s1_1 | _GEN_5366; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9431 = 4'h7 == w_addr_s1_1 | _GEN_5367; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9432 = 4'h8 == w_addr_s1_1 | _GEN_5368; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9433 = 4'h9 == w_addr_s1_1 | _GEN_5369; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9434 = 4'ha == w_addr_s1_1 | _GEN_5370; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9435 = 4'hb == w_addr_s1_1 | _GEN_5371; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9436 = 4'hc == w_addr_s1_1 | _GEN_5372; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9437 = 4'hd == w_addr_s1_1 | _GEN_5373; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9438 = 4'he == w_addr_s1_1 | _GEN_5374; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9439 = 4'hf == w_addr_s1_1 | _GEN_5375; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_339 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_84 = w_valid_s1_1 & _wen_T_339; // @[Sbuffer.scala 156:25]
  wire  _GEN_9488 = 4'h0 == w_addr_s1_1 | _GEN_5424; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9489 = 4'h1 == w_addr_s1_1 | _GEN_5425; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9490 = 4'h2 == w_addr_s1_1 | _GEN_5426; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9491 = 4'h3 == w_addr_s1_1 | _GEN_5427; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9492 = 4'h4 == w_addr_s1_1 | _GEN_5428; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9493 = 4'h5 == w_addr_s1_1 | _GEN_5429; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9494 = 4'h6 == w_addr_s1_1 | _GEN_5430; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9495 = 4'h7 == w_addr_s1_1 | _GEN_5431; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9496 = 4'h8 == w_addr_s1_1 | _GEN_5432; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9497 = 4'h9 == w_addr_s1_1 | _GEN_5433; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9498 = 4'ha == w_addr_s1_1 | _GEN_5434; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9499 = 4'hb == w_addr_s1_1 | _GEN_5435; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9500 = 4'hc == w_addr_s1_1 | _GEN_5436; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9501 = 4'hd == w_addr_s1_1 | _GEN_5437; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9502 = 4'he == w_addr_s1_1 | _GEN_5438; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9503 = 4'hf == w_addr_s1_1 | _GEN_5439; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_343 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_85 = w_valid_s1_1 & _wen_T_343; // @[Sbuffer.scala 156:25]
  wire  _GEN_9552 = 4'h0 == w_addr_s1_1 | _GEN_5488; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9553 = 4'h1 == w_addr_s1_1 | _GEN_5489; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9554 = 4'h2 == w_addr_s1_1 | _GEN_5490; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9555 = 4'h3 == w_addr_s1_1 | _GEN_5491; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9556 = 4'h4 == w_addr_s1_1 | _GEN_5492; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9557 = 4'h5 == w_addr_s1_1 | _GEN_5493; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9558 = 4'h6 == w_addr_s1_1 | _GEN_5494; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9559 = 4'h7 == w_addr_s1_1 | _GEN_5495; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9560 = 4'h8 == w_addr_s1_1 | _GEN_5496; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9561 = 4'h9 == w_addr_s1_1 | _GEN_5497; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9562 = 4'ha == w_addr_s1_1 | _GEN_5498; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9563 = 4'hb == w_addr_s1_1 | _GEN_5499; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9564 = 4'hc == w_addr_s1_1 | _GEN_5500; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9565 = 4'hd == w_addr_s1_1 | _GEN_5501; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9566 = 4'he == w_addr_s1_1 | _GEN_5502; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9567 = 4'hf == w_addr_s1_1 | _GEN_5503; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_347 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_86 = w_valid_s1_1 & _wen_T_347; // @[Sbuffer.scala 156:25]
  wire  _GEN_9616 = 4'h0 == w_addr_s1_1 | _GEN_5552; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9617 = 4'h1 == w_addr_s1_1 | _GEN_5553; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9618 = 4'h2 == w_addr_s1_1 | _GEN_5554; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9619 = 4'h3 == w_addr_s1_1 | _GEN_5555; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9620 = 4'h4 == w_addr_s1_1 | _GEN_5556; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9621 = 4'h5 == w_addr_s1_1 | _GEN_5557; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9622 = 4'h6 == w_addr_s1_1 | _GEN_5558; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9623 = 4'h7 == w_addr_s1_1 | _GEN_5559; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9624 = 4'h8 == w_addr_s1_1 | _GEN_5560; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9625 = 4'h9 == w_addr_s1_1 | _GEN_5561; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9626 = 4'ha == w_addr_s1_1 | _GEN_5562; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9627 = 4'hb == w_addr_s1_1 | _GEN_5563; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9628 = 4'hc == w_addr_s1_1 | _GEN_5564; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9629 = 4'hd == w_addr_s1_1 | _GEN_5565; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9630 = 4'he == w_addr_s1_1 | _GEN_5566; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9631 = 4'hf == w_addr_s1_1 | _GEN_5567; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_351 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h2 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_87 = w_valid_s1_1 & _wen_T_351; // @[Sbuffer.scala 156:25]
  wire  _GEN_9680 = 4'h0 == w_addr_s1_1 | _GEN_5616; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9681 = 4'h1 == w_addr_s1_1 | _GEN_5617; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9682 = 4'h2 == w_addr_s1_1 | _GEN_5618; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9683 = 4'h3 == w_addr_s1_1 | _GEN_5619; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9684 = 4'h4 == w_addr_s1_1 | _GEN_5620; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9685 = 4'h5 == w_addr_s1_1 | _GEN_5621; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9686 = 4'h6 == w_addr_s1_1 | _GEN_5622; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9687 = 4'h7 == w_addr_s1_1 | _GEN_5623; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9688 = 4'h8 == w_addr_s1_1 | _GEN_5624; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9689 = 4'h9 == w_addr_s1_1 | _GEN_5625; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9690 = 4'ha == w_addr_s1_1 | _GEN_5626; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9691 = 4'hb == w_addr_s1_1 | _GEN_5627; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9692 = 4'hc == w_addr_s1_1 | _GEN_5628; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9693 = 4'hd == w_addr_s1_1 | _GEN_5629; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9694 = 4'he == w_addr_s1_1 | _GEN_5630; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9695 = 4'hf == w_addr_s1_1 | _GEN_5631; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_355 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_88 = w_valid_s1_1 & _wen_T_355; // @[Sbuffer.scala 156:25]
  wire  _GEN_9744 = 4'h0 == w_addr_s1_1 | _GEN_5680; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9745 = 4'h1 == w_addr_s1_1 | _GEN_5681; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9746 = 4'h2 == w_addr_s1_1 | _GEN_5682; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9747 = 4'h3 == w_addr_s1_1 | _GEN_5683; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9748 = 4'h4 == w_addr_s1_1 | _GEN_5684; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9749 = 4'h5 == w_addr_s1_1 | _GEN_5685; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9750 = 4'h6 == w_addr_s1_1 | _GEN_5686; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9751 = 4'h7 == w_addr_s1_1 | _GEN_5687; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9752 = 4'h8 == w_addr_s1_1 | _GEN_5688; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9753 = 4'h9 == w_addr_s1_1 | _GEN_5689; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9754 = 4'ha == w_addr_s1_1 | _GEN_5690; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9755 = 4'hb == w_addr_s1_1 | _GEN_5691; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9756 = 4'hc == w_addr_s1_1 | _GEN_5692; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9757 = 4'hd == w_addr_s1_1 | _GEN_5693; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9758 = 4'he == w_addr_s1_1 | _GEN_5694; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9759 = 4'hf == w_addr_s1_1 | _GEN_5695; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_359 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_89 = w_valid_s1_1 & _wen_T_359; // @[Sbuffer.scala 156:25]
  wire  _GEN_9808 = 4'h0 == w_addr_s1_1 | _GEN_5744; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9809 = 4'h1 == w_addr_s1_1 | _GEN_5745; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9810 = 4'h2 == w_addr_s1_1 | _GEN_5746; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9811 = 4'h3 == w_addr_s1_1 | _GEN_5747; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9812 = 4'h4 == w_addr_s1_1 | _GEN_5748; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9813 = 4'h5 == w_addr_s1_1 | _GEN_5749; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9814 = 4'h6 == w_addr_s1_1 | _GEN_5750; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9815 = 4'h7 == w_addr_s1_1 | _GEN_5751; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9816 = 4'h8 == w_addr_s1_1 | _GEN_5752; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9817 = 4'h9 == w_addr_s1_1 | _GEN_5753; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9818 = 4'ha == w_addr_s1_1 | _GEN_5754; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9819 = 4'hb == w_addr_s1_1 | _GEN_5755; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9820 = 4'hc == w_addr_s1_1 | _GEN_5756; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9821 = 4'hd == w_addr_s1_1 | _GEN_5757; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9822 = 4'he == w_addr_s1_1 | _GEN_5758; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9823 = 4'hf == w_addr_s1_1 | _GEN_5759; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_363 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_90 = w_valid_s1_1 & _wen_T_363; // @[Sbuffer.scala 156:25]
  wire  _GEN_9872 = 4'h0 == w_addr_s1_1 | _GEN_5808; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9873 = 4'h1 == w_addr_s1_1 | _GEN_5809; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9874 = 4'h2 == w_addr_s1_1 | _GEN_5810; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9875 = 4'h3 == w_addr_s1_1 | _GEN_5811; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9876 = 4'h4 == w_addr_s1_1 | _GEN_5812; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9877 = 4'h5 == w_addr_s1_1 | _GEN_5813; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9878 = 4'h6 == w_addr_s1_1 | _GEN_5814; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9879 = 4'h7 == w_addr_s1_1 | _GEN_5815; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9880 = 4'h8 == w_addr_s1_1 | _GEN_5816; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9881 = 4'h9 == w_addr_s1_1 | _GEN_5817; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9882 = 4'ha == w_addr_s1_1 | _GEN_5818; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9883 = 4'hb == w_addr_s1_1 | _GEN_5819; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9884 = 4'hc == w_addr_s1_1 | _GEN_5820; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9885 = 4'hd == w_addr_s1_1 | _GEN_5821; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9886 = 4'he == w_addr_s1_1 | _GEN_5822; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9887 = 4'hf == w_addr_s1_1 | _GEN_5823; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_367 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_91 = w_valid_s1_1 & _wen_T_367; // @[Sbuffer.scala 156:25]
  wire  _GEN_9936 = 4'h0 == w_addr_s1_1 | _GEN_5872; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9937 = 4'h1 == w_addr_s1_1 | _GEN_5873; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9938 = 4'h2 == w_addr_s1_1 | _GEN_5874; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9939 = 4'h3 == w_addr_s1_1 | _GEN_5875; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9940 = 4'h4 == w_addr_s1_1 | _GEN_5876; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9941 = 4'h5 == w_addr_s1_1 | _GEN_5877; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9942 = 4'h6 == w_addr_s1_1 | _GEN_5878; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9943 = 4'h7 == w_addr_s1_1 | _GEN_5879; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9944 = 4'h8 == w_addr_s1_1 | _GEN_5880; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9945 = 4'h9 == w_addr_s1_1 | _GEN_5881; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9946 = 4'ha == w_addr_s1_1 | _GEN_5882; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9947 = 4'hb == w_addr_s1_1 | _GEN_5883; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9948 = 4'hc == w_addr_s1_1 | _GEN_5884; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9949 = 4'hd == w_addr_s1_1 | _GEN_5885; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9950 = 4'he == w_addr_s1_1 | _GEN_5886; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_9951 = 4'hf == w_addr_s1_1 | _GEN_5887; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_371 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_92 = w_valid_s1_1 & _wen_T_371; // @[Sbuffer.scala 156:25]
  wire  _GEN_10000 = 4'h0 == w_addr_s1_1 | _GEN_5936; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10001 = 4'h1 == w_addr_s1_1 | _GEN_5937; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10002 = 4'h2 == w_addr_s1_1 | _GEN_5938; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10003 = 4'h3 == w_addr_s1_1 | _GEN_5939; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10004 = 4'h4 == w_addr_s1_1 | _GEN_5940; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10005 = 4'h5 == w_addr_s1_1 | _GEN_5941; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10006 = 4'h6 == w_addr_s1_1 | _GEN_5942; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10007 = 4'h7 == w_addr_s1_1 | _GEN_5943; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10008 = 4'h8 == w_addr_s1_1 | _GEN_5944; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10009 = 4'h9 == w_addr_s1_1 | _GEN_5945; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10010 = 4'ha == w_addr_s1_1 | _GEN_5946; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10011 = 4'hb == w_addr_s1_1 | _GEN_5947; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10012 = 4'hc == w_addr_s1_1 | _GEN_5948; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10013 = 4'hd == w_addr_s1_1 | _GEN_5949; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10014 = 4'he == w_addr_s1_1 | _GEN_5950; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10015 = 4'hf == w_addr_s1_1 | _GEN_5951; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_375 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_93 = w_valid_s1_1 & _wen_T_375; // @[Sbuffer.scala 156:25]
  wire  _GEN_10064 = 4'h0 == w_addr_s1_1 | _GEN_6000; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10065 = 4'h1 == w_addr_s1_1 | _GEN_6001; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10066 = 4'h2 == w_addr_s1_1 | _GEN_6002; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10067 = 4'h3 == w_addr_s1_1 | _GEN_6003; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10068 = 4'h4 == w_addr_s1_1 | _GEN_6004; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10069 = 4'h5 == w_addr_s1_1 | _GEN_6005; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10070 = 4'h6 == w_addr_s1_1 | _GEN_6006; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10071 = 4'h7 == w_addr_s1_1 | _GEN_6007; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10072 = 4'h8 == w_addr_s1_1 | _GEN_6008; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10073 = 4'h9 == w_addr_s1_1 | _GEN_6009; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10074 = 4'ha == w_addr_s1_1 | _GEN_6010; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10075 = 4'hb == w_addr_s1_1 | _GEN_6011; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10076 = 4'hc == w_addr_s1_1 | _GEN_6012; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10077 = 4'hd == w_addr_s1_1 | _GEN_6013; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10078 = 4'he == w_addr_s1_1 | _GEN_6014; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10079 = 4'hf == w_addr_s1_1 | _GEN_6015; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_379 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_94 = w_valid_s1_1 & _wen_T_379; // @[Sbuffer.scala 156:25]
  wire  _GEN_10128 = 4'h0 == w_addr_s1_1 | _GEN_6064; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10129 = 4'h1 == w_addr_s1_1 | _GEN_6065; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10130 = 4'h2 == w_addr_s1_1 | _GEN_6066; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10131 = 4'h3 == w_addr_s1_1 | _GEN_6067; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10132 = 4'h4 == w_addr_s1_1 | _GEN_6068; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10133 = 4'h5 == w_addr_s1_1 | _GEN_6069; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10134 = 4'h6 == w_addr_s1_1 | _GEN_6070; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10135 = 4'h7 == w_addr_s1_1 | _GEN_6071; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10136 = 4'h8 == w_addr_s1_1 | _GEN_6072; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10137 = 4'h9 == w_addr_s1_1 | _GEN_6073; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10138 = 4'ha == w_addr_s1_1 | _GEN_6074; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10139 = 4'hb == w_addr_s1_1 | _GEN_6075; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10140 = 4'hc == w_addr_s1_1 | _GEN_6076; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10141 = 4'hd == w_addr_s1_1 | _GEN_6077; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10142 = 4'he == w_addr_s1_1 | _GEN_6078; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10143 = 4'hf == w_addr_s1_1 | _GEN_6079; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_383 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h3 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_95 = w_valid_s1_1 & _wen_T_383; // @[Sbuffer.scala 156:25]
  wire  _GEN_10192 = 4'h0 == w_addr_s1_1 | _GEN_6128; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10193 = 4'h1 == w_addr_s1_1 | _GEN_6129; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10194 = 4'h2 == w_addr_s1_1 | _GEN_6130; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10195 = 4'h3 == w_addr_s1_1 | _GEN_6131; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10196 = 4'h4 == w_addr_s1_1 | _GEN_6132; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10197 = 4'h5 == w_addr_s1_1 | _GEN_6133; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10198 = 4'h6 == w_addr_s1_1 | _GEN_6134; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10199 = 4'h7 == w_addr_s1_1 | _GEN_6135; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10200 = 4'h8 == w_addr_s1_1 | _GEN_6136; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10201 = 4'h9 == w_addr_s1_1 | _GEN_6137; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10202 = 4'ha == w_addr_s1_1 | _GEN_6138; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10203 = 4'hb == w_addr_s1_1 | _GEN_6139; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10204 = 4'hc == w_addr_s1_1 | _GEN_6140; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10205 = 4'hd == w_addr_s1_1 | _GEN_6141; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10206 = 4'he == w_addr_s1_1 | _GEN_6142; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10207 = 4'hf == w_addr_s1_1 | _GEN_6143; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_387 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_96 = w_valid_s1_1 & _wen_T_387; // @[Sbuffer.scala 156:25]
  wire  _GEN_10256 = 4'h0 == w_addr_s1_1 | _GEN_6192; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10257 = 4'h1 == w_addr_s1_1 | _GEN_6193; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10258 = 4'h2 == w_addr_s1_1 | _GEN_6194; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10259 = 4'h3 == w_addr_s1_1 | _GEN_6195; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10260 = 4'h4 == w_addr_s1_1 | _GEN_6196; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10261 = 4'h5 == w_addr_s1_1 | _GEN_6197; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10262 = 4'h6 == w_addr_s1_1 | _GEN_6198; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10263 = 4'h7 == w_addr_s1_1 | _GEN_6199; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10264 = 4'h8 == w_addr_s1_1 | _GEN_6200; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10265 = 4'h9 == w_addr_s1_1 | _GEN_6201; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10266 = 4'ha == w_addr_s1_1 | _GEN_6202; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10267 = 4'hb == w_addr_s1_1 | _GEN_6203; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10268 = 4'hc == w_addr_s1_1 | _GEN_6204; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10269 = 4'hd == w_addr_s1_1 | _GEN_6205; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10270 = 4'he == w_addr_s1_1 | _GEN_6206; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10271 = 4'hf == w_addr_s1_1 | _GEN_6207; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_391 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_97 = w_valid_s1_1 & _wen_T_391; // @[Sbuffer.scala 156:25]
  wire  _GEN_10320 = 4'h0 == w_addr_s1_1 | _GEN_6256; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10321 = 4'h1 == w_addr_s1_1 | _GEN_6257; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10322 = 4'h2 == w_addr_s1_1 | _GEN_6258; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10323 = 4'h3 == w_addr_s1_1 | _GEN_6259; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10324 = 4'h4 == w_addr_s1_1 | _GEN_6260; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10325 = 4'h5 == w_addr_s1_1 | _GEN_6261; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10326 = 4'h6 == w_addr_s1_1 | _GEN_6262; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10327 = 4'h7 == w_addr_s1_1 | _GEN_6263; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10328 = 4'h8 == w_addr_s1_1 | _GEN_6264; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10329 = 4'h9 == w_addr_s1_1 | _GEN_6265; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10330 = 4'ha == w_addr_s1_1 | _GEN_6266; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10331 = 4'hb == w_addr_s1_1 | _GEN_6267; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10332 = 4'hc == w_addr_s1_1 | _GEN_6268; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10333 = 4'hd == w_addr_s1_1 | _GEN_6269; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10334 = 4'he == w_addr_s1_1 | _GEN_6270; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10335 = 4'hf == w_addr_s1_1 | _GEN_6271; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_395 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_98 = w_valid_s1_1 & _wen_T_395; // @[Sbuffer.scala 156:25]
  wire  _GEN_10384 = 4'h0 == w_addr_s1_1 | _GEN_6320; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10385 = 4'h1 == w_addr_s1_1 | _GEN_6321; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10386 = 4'h2 == w_addr_s1_1 | _GEN_6322; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10387 = 4'h3 == w_addr_s1_1 | _GEN_6323; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10388 = 4'h4 == w_addr_s1_1 | _GEN_6324; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10389 = 4'h5 == w_addr_s1_1 | _GEN_6325; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10390 = 4'h6 == w_addr_s1_1 | _GEN_6326; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10391 = 4'h7 == w_addr_s1_1 | _GEN_6327; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10392 = 4'h8 == w_addr_s1_1 | _GEN_6328; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10393 = 4'h9 == w_addr_s1_1 | _GEN_6329; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10394 = 4'ha == w_addr_s1_1 | _GEN_6330; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10395 = 4'hb == w_addr_s1_1 | _GEN_6331; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10396 = 4'hc == w_addr_s1_1 | _GEN_6332; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10397 = 4'hd == w_addr_s1_1 | _GEN_6333; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10398 = 4'he == w_addr_s1_1 | _GEN_6334; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10399 = 4'hf == w_addr_s1_1 | _GEN_6335; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_399 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_99 = w_valid_s1_1 & _wen_T_399; // @[Sbuffer.scala 156:25]
  wire  _GEN_10448 = 4'h0 == w_addr_s1_1 | _GEN_6384; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10449 = 4'h1 == w_addr_s1_1 | _GEN_6385; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10450 = 4'h2 == w_addr_s1_1 | _GEN_6386; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10451 = 4'h3 == w_addr_s1_1 | _GEN_6387; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10452 = 4'h4 == w_addr_s1_1 | _GEN_6388; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10453 = 4'h5 == w_addr_s1_1 | _GEN_6389; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10454 = 4'h6 == w_addr_s1_1 | _GEN_6390; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10455 = 4'h7 == w_addr_s1_1 | _GEN_6391; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10456 = 4'h8 == w_addr_s1_1 | _GEN_6392; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10457 = 4'h9 == w_addr_s1_1 | _GEN_6393; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10458 = 4'ha == w_addr_s1_1 | _GEN_6394; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10459 = 4'hb == w_addr_s1_1 | _GEN_6395; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10460 = 4'hc == w_addr_s1_1 | _GEN_6396; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10461 = 4'hd == w_addr_s1_1 | _GEN_6397; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10462 = 4'he == w_addr_s1_1 | _GEN_6398; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10463 = 4'hf == w_addr_s1_1 | _GEN_6399; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_403 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_100 = w_valid_s1_1 & _wen_T_403; // @[Sbuffer.scala 156:25]
  wire  _GEN_10512 = 4'h0 == w_addr_s1_1 | _GEN_6448; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10513 = 4'h1 == w_addr_s1_1 | _GEN_6449; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10514 = 4'h2 == w_addr_s1_1 | _GEN_6450; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10515 = 4'h3 == w_addr_s1_1 | _GEN_6451; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10516 = 4'h4 == w_addr_s1_1 | _GEN_6452; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10517 = 4'h5 == w_addr_s1_1 | _GEN_6453; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10518 = 4'h6 == w_addr_s1_1 | _GEN_6454; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10519 = 4'h7 == w_addr_s1_1 | _GEN_6455; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10520 = 4'h8 == w_addr_s1_1 | _GEN_6456; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10521 = 4'h9 == w_addr_s1_1 | _GEN_6457; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10522 = 4'ha == w_addr_s1_1 | _GEN_6458; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10523 = 4'hb == w_addr_s1_1 | _GEN_6459; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10524 = 4'hc == w_addr_s1_1 | _GEN_6460; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10525 = 4'hd == w_addr_s1_1 | _GEN_6461; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10526 = 4'he == w_addr_s1_1 | _GEN_6462; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10527 = 4'hf == w_addr_s1_1 | _GEN_6463; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_407 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_101 = w_valid_s1_1 & _wen_T_407; // @[Sbuffer.scala 156:25]
  wire  _GEN_10576 = 4'h0 == w_addr_s1_1 | _GEN_6512; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10577 = 4'h1 == w_addr_s1_1 | _GEN_6513; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10578 = 4'h2 == w_addr_s1_1 | _GEN_6514; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10579 = 4'h3 == w_addr_s1_1 | _GEN_6515; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10580 = 4'h4 == w_addr_s1_1 | _GEN_6516; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10581 = 4'h5 == w_addr_s1_1 | _GEN_6517; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10582 = 4'h6 == w_addr_s1_1 | _GEN_6518; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10583 = 4'h7 == w_addr_s1_1 | _GEN_6519; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10584 = 4'h8 == w_addr_s1_1 | _GEN_6520; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10585 = 4'h9 == w_addr_s1_1 | _GEN_6521; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10586 = 4'ha == w_addr_s1_1 | _GEN_6522; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10587 = 4'hb == w_addr_s1_1 | _GEN_6523; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10588 = 4'hc == w_addr_s1_1 | _GEN_6524; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10589 = 4'hd == w_addr_s1_1 | _GEN_6525; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10590 = 4'he == w_addr_s1_1 | _GEN_6526; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10591 = 4'hf == w_addr_s1_1 | _GEN_6527; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_411 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_102 = w_valid_s1_1 & _wen_T_411; // @[Sbuffer.scala 156:25]
  wire  _GEN_10640 = 4'h0 == w_addr_s1_1 | _GEN_6576; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10641 = 4'h1 == w_addr_s1_1 | _GEN_6577; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10642 = 4'h2 == w_addr_s1_1 | _GEN_6578; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10643 = 4'h3 == w_addr_s1_1 | _GEN_6579; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10644 = 4'h4 == w_addr_s1_1 | _GEN_6580; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10645 = 4'h5 == w_addr_s1_1 | _GEN_6581; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10646 = 4'h6 == w_addr_s1_1 | _GEN_6582; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10647 = 4'h7 == w_addr_s1_1 | _GEN_6583; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10648 = 4'h8 == w_addr_s1_1 | _GEN_6584; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10649 = 4'h9 == w_addr_s1_1 | _GEN_6585; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10650 = 4'ha == w_addr_s1_1 | _GEN_6586; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10651 = 4'hb == w_addr_s1_1 | _GEN_6587; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10652 = 4'hc == w_addr_s1_1 | _GEN_6588; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10653 = 4'hd == w_addr_s1_1 | _GEN_6589; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10654 = 4'he == w_addr_s1_1 | _GEN_6590; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10655 = 4'hf == w_addr_s1_1 | _GEN_6591; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_415 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h4 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_103 = w_valid_s1_1 & _wen_T_415; // @[Sbuffer.scala 156:25]
  wire  _GEN_10704 = 4'h0 == w_addr_s1_1 | _GEN_6640; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10705 = 4'h1 == w_addr_s1_1 | _GEN_6641; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10706 = 4'h2 == w_addr_s1_1 | _GEN_6642; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10707 = 4'h3 == w_addr_s1_1 | _GEN_6643; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10708 = 4'h4 == w_addr_s1_1 | _GEN_6644; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10709 = 4'h5 == w_addr_s1_1 | _GEN_6645; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10710 = 4'h6 == w_addr_s1_1 | _GEN_6646; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10711 = 4'h7 == w_addr_s1_1 | _GEN_6647; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10712 = 4'h8 == w_addr_s1_1 | _GEN_6648; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10713 = 4'h9 == w_addr_s1_1 | _GEN_6649; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10714 = 4'ha == w_addr_s1_1 | _GEN_6650; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10715 = 4'hb == w_addr_s1_1 | _GEN_6651; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10716 = 4'hc == w_addr_s1_1 | _GEN_6652; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10717 = 4'hd == w_addr_s1_1 | _GEN_6653; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10718 = 4'he == w_addr_s1_1 | _GEN_6654; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10719 = 4'hf == w_addr_s1_1 | _GEN_6655; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_419 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_104 = w_valid_s1_1 & _wen_T_419; // @[Sbuffer.scala 156:25]
  wire  _GEN_10768 = 4'h0 == w_addr_s1_1 | _GEN_6704; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10769 = 4'h1 == w_addr_s1_1 | _GEN_6705; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10770 = 4'h2 == w_addr_s1_1 | _GEN_6706; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10771 = 4'h3 == w_addr_s1_1 | _GEN_6707; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10772 = 4'h4 == w_addr_s1_1 | _GEN_6708; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10773 = 4'h5 == w_addr_s1_1 | _GEN_6709; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10774 = 4'h6 == w_addr_s1_1 | _GEN_6710; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10775 = 4'h7 == w_addr_s1_1 | _GEN_6711; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10776 = 4'h8 == w_addr_s1_1 | _GEN_6712; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10777 = 4'h9 == w_addr_s1_1 | _GEN_6713; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10778 = 4'ha == w_addr_s1_1 | _GEN_6714; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10779 = 4'hb == w_addr_s1_1 | _GEN_6715; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10780 = 4'hc == w_addr_s1_1 | _GEN_6716; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10781 = 4'hd == w_addr_s1_1 | _GEN_6717; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10782 = 4'he == w_addr_s1_1 | _GEN_6718; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10783 = 4'hf == w_addr_s1_1 | _GEN_6719; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_423 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_105 = w_valid_s1_1 & _wen_T_423; // @[Sbuffer.scala 156:25]
  wire  _GEN_10832 = 4'h0 == w_addr_s1_1 | _GEN_6768; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10833 = 4'h1 == w_addr_s1_1 | _GEN_6769; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10834 = 4'h2 == w_addr_s1_1 | _GEN_6770; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10835 = 4'h3 == w_addr_s1_1 | _GEN_6771; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10836 = 4'h4 == w_addr_s1_1 | _GEN_6772; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10837 = 4'h5 == w_addr_s1_1 | _GEN_6773; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10838 = 4'h6 == w_addr_s1_1 | _GEN_6774; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10839 = 4'h7 == w_addr_s1_1 | _GEN_6775; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10840 = 4'h8 == w_addr_s1_1 | _GEN_6776; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10841 = 4'h9 == w_addr_s1_1 | _GEN_6777; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10842 = 4'ha == w_addr_s1_1 | _GEN_6778; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10843 = 4'hb == w_addr_s1_1 | _GEN_6779; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10844 = 4'hc == w_addr_s1_1 | _GEN_6780; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10845 = 4'hd == w_addr_s1_1 | _GEN_6781; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10846 = 4'he == w_addr_s1_1 | _GEN_6782; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10847 = 4'hf == w_addr_s1_1 | _GEN_6783; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_427 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_106 = w_valid_s1_1 & _wen_T_427; // @[Sbuffer.scala 156:25]
  wire  _GEN_10896 = 4'h0 == w_addr_s1_1 | _GEN_6832; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10897 = 4'h1 == w_addr_s1_1 | _GEN_6833; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10898 = 4'h2 == w_addr_s1_1 | _GEN_6834; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10899 = 4'h3 == w_addr_s1_1 | _GEN_6835; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10900 = 4'h4 == w_addr_s1_1 | _GEN_6836; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10901 = 4'h5 == w_addr_s1_1 | _GEN_6837; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10902 = 4'h6 == w_addr_s1_1 | _GEN_6838; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10903 = 4'h7 == w_addr_s1_1 | _GEN_6839; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10904 = 4'h8 == w_addr_s1_1 | _GEN_6840; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10905 = 4'h9 == w_addr_s1_1 | _GEN_6841; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10906 = 4'ha == w_addr_s1_1 | _GEN_6842; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10907 = 4'hb == w_addr_s1_1 | _GEN_6843; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10908 = 4'hc == w_addr_s1_1 | _GEN_6844; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10909 = 4'hd == w_addr_s1_1 | _GEN_6845; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10910 = 4'he == w_addr_s1_1 | _GEN_6846; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10911 = 4'hf == w_addr_s1_1 | _GEN_6847; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_431 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_107 = w_valid_s1_1 & _wen_T_431; // @[Sbuffer.scala 156:25]
  wire  _GEN_10960 = 4'h0 == w_addr_s1_1 | _GEN_6896; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10961 = 4'h1 == w_addr_s1_1 | _GEN_6897; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10962 = 4'h2 == w_addr_s1_1 | _GEN_6898; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10963 = 4'h3 == w_addr_s1_1 | _GEN_6899; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10964 = 4'h4 == w_addr_s1_1 | _GEN_6900; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10965 = 4'h5 == w_addr_s1_1 | _GEN_6901; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10966 = 4'h6 == w_addr_s1_1 | _GEN_6902; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10967 = 4'h7 == w_addr_s1_1 | _GEN_6903; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10968 = 4'h8 == w_addr_s1_1 | _GEN_6904; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10969 = 4'h9 == w_addr_s1_1 | _GEN_6905; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10970 = 4'ha == w_addr_s1_1 | _GEN_6906; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10971 = 4'hb == w_addr_s1_1 | _GEN_6907; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10972 = 4'hc == w_addr_s1_1 | _GEN_6908; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10973 = 4'hd == w_addr_s1_1 | _GEN_6909; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10974 = 4'he == w_addr_s1_1 | _GEN_6910; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_10975 = 4'hf == w_addr_s1_1 | _GEN_6911; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_435 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_108 = w_valid_s1_1 & _wen_T_435; // @[Sbuffer.scala 156:25]
  wire  _GEN_11024 = 4'h0 == w_addr_s1_1 | _GEN_6960; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11025 = 4'h1 == w_addr_s1_1 | _GEN_6961; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11026 = 4'h2 == w_addr_s1_1 | _GEN_6962; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11027 = 4'h3 == w_addr_s1_1 | _GEN_6963; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11028 = 4'h4 == w_addr_s1_1 | _GEN_6964; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11029 = 4'h5 == w_addr_s1_1 | _GEN_6965; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11030 = 4'h6 == w_addr_s1_1 | _GEN_6966; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11031 = 4'h7 == w_addr_s1_1 | _GEN_6967; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11032 = 4'h8 == w_addr_s1_1 | _GEN_6968; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11033 = 4'h9 == w_addr_s1_1 | _GEN_6969; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11034 = 4'ha == w_addr_s1_1 | _GEN_6970; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11035 = 4'hb == w_addr_s1_1 | _GEN_6971; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11036 = 4'hc == w_addr_s1_1 | _GEN_6972; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11037 = 4'hd == w_addr_s1_1 | _GEN_6973; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11038 = 4'he == w_addr_s1_1 | _GEN_6974; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11039 = 4'hf == w_addr_s1_1 | _GEN_6975; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_439 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_109 = w_valid_s1_1 & _wen_T_439; // @[Sbuffer.scala 156:25]
  wire  _GEN_11088 = 4'h0 == w_addr_s1_1 | _GEN_7024; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11089 = 4'h1 == w_addr_s1_1 | _GEN_7025; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11090 = 4'h2 == w_addr_s1_1 | _GEN_7026; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11091 = 4'h3 == w_addr_s1_1 | _GEN_7027; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11092 = 4'h4 == w_addr_s1_1 | _GEN_7028; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11093 = 4'h5 == w_addr_s1_1 | _GEN_7029; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11094 = 4'h6 == w_addr_s1_1 | _GEN_7030; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11095 = 4'h7 == w_addr_s1_1 | _GEN_7031; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11096 = 4'h8 == w_addr_s1_1 | _GEN_7032; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11097 = 4'h9 == w_addr_s1_1 | _GEN_7033; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11098 = 4'ha == w_addr_s1_1 | _GEN_7034; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11099 = 4'hb == w_addr_s1_1 | _GEN_7035; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11100 = 4'hc == w_addr_s1_1 | _GEN_7036; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11101 = 4'hd == w_addr_s1_1 | _GEN_7037; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11102 = 4'he == w_addr_s1_1 | _GEN_7038; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11103 = 4'hf == w_addr_s1_1 | _GEN_7039; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_443 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_110 = w_valid_s1_1 & _wen_T_443; // @[Sbuffer.scala 156:25]
  wire  _GEN_11152 = 4'h0 == w_addr_s1_1 | _GEN_7088; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11153 = 4'h1 == w_addr_s1_1 | _GEN_7089; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11154 = 4'h2 == w_addr_s1_1 | _GEN_7090; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11155 = 4'h3 == w_addr_s1_1 | _GEN_7091; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11156 = 4'h4 == w_addr_s1_1 | _GEN_7092; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11157 = 4'h5 == w_addr_s1_1 | _GEN_7093; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11158 = 4'h6 == w_addr_s1_1 | _GEN_7094; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11159 = 4'h7 == w_addr_s1_1 | _GEN_7095; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11160 = 4'h8 == w_addr_s1_1 | _GEN_7096; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11161 = 4'h9 == w_addr_s1_1 | _GEN_7097; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11162 = 4'ha == w_addr_s1_1 | _GEN_7098; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11163 = 4'hb == w_addr_s1_1 | _GEN_7099; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11164 = 4'hc == w_addr_s1_1 | _GEN_7100; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11165 = 4'hd == w_addr_s1_1 | _GEN_7101; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11166 = 4'he == w_addr_s1_1 | _GEN_7102; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11167 = 4'hf == w_addr_s1_1 | _GEN_7103; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_447 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h5 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_111 = w_valid_s1_1 & _wen_T_447; // @[Sbuffer.scala 156:25]
  wire  _GEN_11216 = 4'h0 == w_addr_s1_1 | _GEN_7152; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11217 = 4'h1 == w_addr_s1_1 | _GEN_7153; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11218 = 4'h2 == w_addr_s1_1 | _GEN_7154; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11219 = 4'h3 == w_addr_s1_1 | _GEN_7155; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11220 = 4'h4 == w_addr_s1_1 | _GEN_7156; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11221 = 4'h5 == w_addr_s1_1 | _GEN_7157; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11222 = 4'h6 == w_addr_s1_1 | _GEN_7158; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11223 = 4'h7 == w_addr_s1_1 | _GEN_7159; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11224 = 4'h8 == w_addr_s1_1 | _GEN_7160; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11225 = 4'h9 == w_addr_s1_1 | _GEN_7161; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11226 = 4'ha == w_addr_s1_1 | _GEN_7162; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11227 = 4'hb == w_addr_s1_1 | _GEN_7163; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11228 = 4'hc == w_addr_s1_1 | _GEN_7164; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11229 = 4'hd == w_addr_s1_1 | _GEN_7165; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11230 = 4'he == w_addr_s1_1 | _GEN_7166; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11231 = 4'hf == w_addr_s1_1 | _GEN_7167; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_451 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_112 = w_valid_s1_1 & _wen_T_451; // @[Sbuffer.scala 156:25]
  wire  _GEN_11280 = 4'h0 == w_addr_s1_1 | _GEN_7216; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11281 = 4'h1 == w_addr_s1_1 | _GEN_7217; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11282 = 4'h2 == w_addr_s1_1 | _GEN_7218; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11283 = 4'h3 == w_addr_s1_1 | _GEN_7219; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11284 = 4'h4 == w_addr_s1_1 | _GEN_7220; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11285 = 4'h5 == w_addr_s1_1 | _GEN_7221; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11286 = 4'h6 == w_addr_s1_1 | _GEN_7222; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11287 = 4'h7 == w_addr_s1_1 | _GEN_7223; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11288 = 4'h8 == w_addr_s1_1 | _GEN_7224; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11289 = 4'h9 == w_addr_s1_1 | _GEN_7225; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11290 = 4'ha == w_addr_s1_1 | _GEN_7226; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11291 = 4'hb == w_addr_s1_1 | _GEN_7227; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11292 = 4'hc == w_addr_s1_1 | _GEN_7228; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11293 = 4'hd == w_addr_s1_1 | _GEN_7229; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11294 = 4'he == w_addr_s1_1 | _GEN_7230; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11295 = 4'hf == w_addr_s1_1 | _GEN_7231; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_455 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_113 = w_valid_s1_1 & _wen_T_455; // @[Sbuffer.scala 156:25]
  wire  _GEN_11344 = 4'h0 == w_addr_s1_1 | _GEN_7280; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11345 = 4'h1 == w_addr_s1_1 | _GEN_7281; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11346 = 4'h2 == w_addr_s1_1 | _GEN_7282; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11347 = 4'h3 == w_addr_s1_1 | _GEN_7283; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11348 = 4'h4 == w_addr_s1_1 | _GEN_7284; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11349 = 4'h5 == w_addr_s1_1 | _GEN_7285; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11350 = 4'h6 == w_addr_s1_1 | _GEN_7286; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11351 = 4'h7 == w_addr_s1_1 | _GEN_7287; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11352 = 4'h8 == w_addr_s1_1 | _GEN_7288; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11353 = 4'h9 == w_addr_s1_1 | _GEN_7289; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11354 = 4'ha == w_addr_s1_1 | _GEN_7290; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11355 = 4'hb == w_addr_s1_1 | _GEN_7291; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11356 = 4'hc == w_addr_s1_1 | _GEN_7292; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11357 = 4'hd == w_addr_s1_1 | _GEN_7293; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11358 = 4'he == w_addr_s1_1 | _GEN_7294; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11359 = 4'hf == w_addr_s1_1 | _GEN_7295; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_459 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_114 = w_valid_s1_1 & _wen_T_459; // @[Sbuffer.scala 156:25]
  wire  _GEN_11408 = 4'h0 == w_addr_s1_1 | _GEN_7344; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11409 = 4'h1 == w_addr_s1_1 | _GEN_7345; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11410 = 4'h2 == w_addr_s1_1 | _GEN_7346; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11411 = 4'h3 == w_addr_s1_1 | _GEN_7347; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11412 = 4'h4 == w_addr_s1_1 | _GEN_7348; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11413 = 4'h5 == w_addr_s1_1 | _GEN_7349; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11414 = 4'h6 == w_addr_s1_1 | _GEN_7350; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11415 = 4'h7 == w_addr_s1_1 | _GEN_7351; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11416 = 4'h8 == w_addr_s1_1 | _GEN_7352; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11417 = 4'h9 == w_addr_s1_1 | _GEN_7353; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11418 = 4'ha == w_addr_s1_1 | _GEN_7354; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11419 = 4'hb == w_addr_s1_1 | _GEN_7355; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11420 = 4'hc == w_addr_s1_1 | _GEN_7356; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11421 = 4'hd == w_addr_s1_1 | _GEN_7357; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11422 = 4'he == w_addr_s1_1 | _GEN_7358; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11423 = 4'hf == w_addr_s1_1 | _GEN_7359; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_463 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_115 = w_valid_s1_1 & _wen_T_463; // @[Sbuffer.scala 156:25]
  wire  _GEN_11472 = 4'h0 == w_addr_s1_1 | _GEN_7408; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11473 = 4'h1 == w_addr_s1_1 | _GEN_7409; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11474 = 4'h2 == w_addr_s1_1 | _GEN_7410; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11475 = 4'h3 == w_addr_s1_1 | _GEN_7411; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11476 = 4'h4 == w_addr_s1_1 | _GEN_7412; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11477 = 4'h5 == w_addr_s1_1 | _GEN_7413; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11478 = 4'h6 == w_addr_s1_1 | _GEN_7414; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11479 = 4'h7 == w_addr_s1_1 | _GEN_7415; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11480 = 4'h8 == w_addr_s1_1 | _GEN_7416; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11481 = 4'h9 == w_addr_s1_1 | _GEN_7417; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11482 = 4'ha == w_addr_s1_1 | _GEN_7418; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11483 = 4'hb == w_addr_s1_1 | _GEN_7419; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11484 = 4'hc == w_addr_s1_1 | _GEN_7420; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11485 = 4'hd == w_addr_s1_1 | _GEN_7421; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11486 = 4'he == w_addr_s1_1 | _GEN_7422; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11487 = 4'hf == w_addr_s1_1 | _GEN_7423; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_467 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_116 = w_valid_s1_1 & _wen_T_467; // @[Sbuffer.scala 156:25]
  wire  _GEN_11536 = 4'h0 == w_addr_s1_1 | _GEN_7472; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11537 = 4'h1 == w_addr_s1_1 | _GEN_7473; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11538 = 4'h2 == w_addr_s1_1 | _GEN_7474; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11539 = 4'h3 == w_addr_s1_1 | _GEN_7475; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11540 = 4'h4 == w_addr_s1_1 | _GEN_7476; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11541 = 4'h5 == w_addr_s1_1 | _GEN_7477; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11542 = 4'h6 == w_addr_s1_1 | _GEN_7478; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11543 = 4'h7 == w_addr_s1_1 | _GEN_7479; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11544 = 4'h8 == w_addr_s1_1 | _GEN_7480; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11545 = 4'h9 == w_addr_s1_1 | _GEN_7481; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11546 = 4'ha == w_addr_s1_1 | _GEN_7482; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11547 = 4'hb == w_addr_s1_1 | _GEN_7483; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11548 = 4'hc == w_addr_s1_1 | _GEN_7484; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11549 = 4'hd == w_addr_s1_1 | _GEN_7485; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11550 = 4'he == w_addr_s1_1 | _GEN_7486; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11551 = 4'hf == w_addr_s1_1 | _GEN_7487; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_471 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_117 = w_valid_s1_1 & _wen_T_471; // @[Sbuffer.scala 156:25]
  wire  _GEN_11600 = 4'h0 == w_addr_s1_1 | _GEN_7536; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11601 = 4'h1 == w_addr_s1_1 | _GEN_7537; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11602 = 4'h2 == w_addr_s1_1 | _GEN_7538; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11603 = 4'h3 == w_addr_s1_1 | _GEN_7539; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11604 = 4'h4 == w_addr_s1_1 | _GEN_7540; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11605 = 4'h5 == w_addr_s1_1 | _GEN_7541; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11606 = 4'h6 == w_addr_s1_1 | _GEN_7542; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11607 = 4'h7 == w_addr_s1_1 | _GEN_7543; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11608 = 4'h8 == w_addr_s1_1 | _GEN_7544; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11609 = 4'h9 == w_addr_s1_1 | _GEN_7545; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11610 = 4'ha == w_addr_s1_1 | _GEN_7546; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11611 = 4'hb == w_addr_s1_1 | _GEN_7547; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11612 = 4'hc == w_addr_s1_1 | _GEN_7548; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11613 = 4'hd == w_addr_s1_1 | _GEN_7549; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11614 = 4'he == w_addr_s1_1 | _GEN_7550; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11615 = 4'hf == w_addr_s1_1 | _GEN_7551; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_475 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_118 = w_valid_s1_1 & _wen_T_475; // @[Sbuffer.scala 156:25]
  wire  _GEN_11664 = 4'h0 == w_addr_s1_1 | _GEN_7600; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11665 = 4'h1 == w_addr_s1_1 | _GEN_7601; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11666 = 4'h2 == w_addr_s1_1 | _GEN_7602; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11667 = 4'h3 == w_addr_s1_1 | _GEN_7603; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11668 = 4'h4 == w_addr_s1_1 | _GEN_7604; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11669 = 4'h5 == w_addr_s1_1 | _GEN_7605; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11670 = 4'h6 == w_addr_s1_1 | _GEN_7606; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11671 = 4'h7 == w_addr_s1_1 | _GEN_7607; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11672 = 4'h8 == w_addr_s1_1 | _GEN_7608; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11673 = 4'h9 == w_addr_s1_1 | _GEN_7609; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11674 = 4'ha == w_addr_s1_1 | _GEN_7610; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11675 = 4'hb == w_addr_s1_1 | _GEN_7611; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11676 = 4'hc == w_addr_s1_1 | _GEN_7612; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11677 = 4'hd == w_addr_s1_1 | _GEN_7613; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11678 = 4'he == w_addr_s1_1 | _GEN_7614; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11679 = 4'hf == w_addr_s1_1 | _GEN_7615; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_479 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h6 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_119 = w_valid_s1_1 & _wen_T_479; // @[Sbuffer.scala 156:25]
  wire  _GEN_11728 = 4'h0 == w_addr_s1_1 | _GEN_7664; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11729 = 4'h1 == w_addr_s1_1 | _GEN_7665; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11730 = 4'h2 == w_addr_s1_1 | _GEN_7666; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11731 = 4'h3 == w_addr_s1_1 | _GEN_7667; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11732 = 4'h4 == w_addr_s1_1 | _GEN_7668; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11733 = 4'h5 == w_addr_s1_1 | _GEN_7669; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11734 = 4'h6 == w_addr_s1_1 | _GEN_7670; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11735 = 4'h7 == w_addr_s1_1 | _GEN_7671; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11736 = 4'h8 == w_addr_s1_1 | _GEN_7672; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11737 = 4'h9 == w_addr_s1_1 | _GEN_7673; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11738 = 4'ha == w_addr_s1_1 | _GEN_7674; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11739 = 4'hb == w_addr_s1_1 | _GEN_7675; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11740 = 4'hc == w_addr_s1_1 | _GEN_7676; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11741 = 4'hd == w_addr_s1_1 | _GEN_7677; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11742 = 4'he == w_addr_s1_1 | _GEN_7678; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11743 = 4'hf == w_addr_s1_1 | _GEN_7679; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_483 = w_mask_s1_1[0] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_120 = w_valid_s1_1 & _wen_T_483; // @[Sbuffer.scala 156:25]
  wire  _GEN_11792 = 4'h0 == w_addr_s1_1 | _GEN_7728; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11793 = 4'h1 == w_addr_s1_1 | _GEN_7729; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11794 = 4'h2 == w_addr_s1_1 | _GEN_7730; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11795 = 4'h3 == w_addr_s1_1 | _GEN_7731; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11796 = 4'h4 == w_addr_s1_1 | _GEN_7732; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11797 = 4'h5 == w_addr_s1_1 | _GEN_7733; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11798 = 4'h6 == w_addr_s1_1 | _GEN_7734; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11799 = 4'h7 == w_addr_s1_1 | _GEN_7735; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11800 = 4'h8 == w_addr_s1_1 | _GEN_7736; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11801 = 4'h9 == w_addr_s1_1 | _GEN_7737; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11802 = 4'ha == w_addr_s1_1 | _GEN_7738; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11803 = 4'hb == w_addr_s1_1 | _GEN_7739; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11804 = 4'hc == w_addr_s1_1 | _GEN_7740; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11805 = 4'hd == w_addr_s1_1 | _GEN_7741; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11806 = 4'he == w_addr_s1_1 | _GEN_7742; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11807 = 4'hf == w_addr_s1_1 | _GEN_7743; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_487 = w_mask_s1_1[1] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_121 = w_valid_s1_1 & _wen_T_487; // @[Sbuffer.scala 156:25]
  wire  _GEN_11856 = 4'h0 == w_addr_s1_1 | _GEN_7792; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11857 = 4'h1 == w_addr_s1_1 | _GEN_7793; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11858 = 4'h2 == w_addr_s1_1 | _GEN_7794; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11859 = 4'h3 == w_addr_s1_1 | _GEN_7795; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11860 = 4'h4 == w_addr_s1_1 | _GEN_7796; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11861 = 4'h5 == w_addr_s1_1 | _GEN_7797; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11862 = 4'h6 == w_addr_s1_1 | _GEN_7798; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11863 = 4'h7 == w_addr_s1_1 | _GEN_7799; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11864 = 4'h8 == w_addr_s1_1 | _GEN_7800; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11865 = 4'h9 == w_addr_s1_1 | _GEN_7801; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11866 = 4'ha == w_addr_s1_1 | _GEN_7802; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11867 = 4'hb == w_addr_s1_1 | _GEN_7803; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11868 = 4'hc == w_addr_s1_1 | _GEN_7804; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11869 = 4'hd == w_addr_s1_1 | _GEN_7805; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11870 = 4'he == w_addr_s1_1 | _GEN_7806; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11871 = 4'hf == w_addr_s1_1 | _GEN_7807; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_491 = w_mask_s1_1[2] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_122 = w_valid_s1_1 & _wen_T_491; // @[Sbuffer.scala 156:25]
  wire  _GEN_11920 = 4'h0 == w_addr_s1_1 | _GEN_7856; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11921 = 4'h1 == w_addr_s1_1 | _GEN_7857; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11922 = 4'h2 == w_addr_s1_1 | _GEN_7858; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11923 = 4'h3 == w_addr_s1_1 | _GEN_7859; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11924 = 4'h4 == w_addr_s1_1 | _GEN_7860; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11925 = 4'h5 == w_addr_s1_1 | _GEN_7861; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11926 = 4'h6 == w_addr_s1_1 | _GEN_7862; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11927 = 4'h7 == w_addr_s1_1 | _GEN_7863; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11928 = 4'h8 == w_addr_s1_1 | _GEN_7864; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11929 = 4'h9 == w_addr_s1_1 | _GEN_7865; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11930 = 4'ha == w_addr_s1_1 | _GEN_7866; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11931 = 4'hb == w_addr_s1_1 | _GEN_7867; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11932 = 4'hc == w_addr_s1_1 | _GEN_7868; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11933 = 4'hd == w_addr_s1_1 | _GEN_7869; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11934 = 4'he == w_addr_s1_1 | _GEN_7870; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11935 = 4'hf == w_addr_s1_1 | _GEN_7871; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_495 = w_mask_s1_1[3] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_123 = w_valid_s1_1 & _wen_T_495; // @[Sbuffer.scala 156:25]
  wire  _GEN_11984 = 4'h0 == w_addr_s1_1 | _GEN_7920; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11985 = 4'h1 == w_addr_s1_1 | _GEN_7921; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11986 = 4'h2 == w_addr_s1_1 | _GEN_7922; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11987 = 4'h3 == w_addr_s1_1 | _GEN_7923; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11988 = 4'h4 == w_addr_s1_1 | _GEN_7924; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11989 = 4'h5 == w_addr_s1_1 | _GEN_7925; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11990 = 4'h6 == w_addr_s1_1 | _GEN_7926; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11991 = 4'h7 == w_addr_s1_1 | _GEN_7927; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11992 = 4'h8 == w_addr_s1_1 | _GEN_7928; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11993 = 4'h9 == w_addr_s1_1 | _GEN_7929; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11994 = 4'ha == w_addr_s1_1 | _GEN_7930; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11995 = 4'hb == w_addr_s1_1 | _GEN_7931; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11996 = 4'hc == w_addr_s1_1 | _GEN_7932; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11997 = 4'hd == w_addr_s1_1 | _GEN_7933; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11998 = 4'he == w_addr_s1_1 | _GEN_7934; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_11999 = 4'hf == w_addr_s1_1 | _GEN_7935; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_499 = w_mask_s1_1[4] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_124 = w_valid_s1_1 & _wen_T_499; // @[Sbuffer.scala 156:25]
  wire  _GEN_12048 = 4'h0 == w_addr_s1_1 | _GEN_7984; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12049 = 4'h1 == w_addr_s1_1 | _GEN_7985; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12050 = 4'h2 == w_addr_s1_1 | _GEN_7986; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12051 = 4'h3 == w_addr_s1_1 | _GEN_7987; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12052 = 4'h4 == w_addr_s1_1 | _GEN_7988; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12053 = 4'h5 == w_addr_s1_1 | _GEN_7989; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12054 = 4'h6 == w_addr_s1_1 | _GEN_7990; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12055 = 4'h7 == w_addr_s1_1 | _GEN_7991; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12056 = 4'h8 == w_addr_s1_1 | _GEN_7992; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12057 = 4'h9 == w_addr_s1_1 | _GEN_7993; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12058 = 4'ha == w_addr_s1_1 | _GEN_7994; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12059 = 4'hb == w_addr_s1_1 | _GEN_7995; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12060 = 4'hc == w_addr_s1_1 | _GEN_7996; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12061 = 4'hd == w_addr_s1_1 | _GEN_7997; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12062 = 4'he == w_addr_s1_1 | _GEN_7998; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12063 = 4'hf == w_addr_s1_1 | _GEN_7999; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_503 = w_mask_s1_1[5] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_125 = w_valid_s1_1 & _wen_T_503; // @[Sbuffer.scala 156:25]
  wire  _GEN_12112 = 4'h0 == w_addr_s1_1 | _GEN_8048; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12113 = 4'h1 == w_addr_s1_1 | _GEN_8049; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12114 = 4'h2 == w_addr_s1_1 | _GEN_8050; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12115 = 4'h3 == w_addr_s1_1 | _GEN_8051; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12116 = 4'h4 == w_addr_s1_1 | _GEN_8052; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12117 = 4'h5 == w_addr_s1_1 | _GEN_8053; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12118 = 4'h6 == w_addr_s1_1 | _GEN_8054; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12119 = 4'h7 == w_addr_s1_1 | _GEN_8055; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12120 = 4'h8 == w_addr_s1_1 | _GEN_8056; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12121 = 4'h9 == w_addr_s1_1 | _GEN_8057; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12122 = 4'ha == w_addr_s1_1 | _GEN_8058; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12123 = 4'hb == w_addr_s1_1 | _GEN_8059; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12124 = 4'hc == w_addr_s1_1 | _GEN_8060; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12125 = 4'hd == w_addr_s1_1 | _GEN_8061; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12126 = 4'he == w_addr_s1_1 | _GEN_8062; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12127 = 4'hf == w_addr_s1_1 | _GEN_8063; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_507 = w_mask_s1_1[6] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_126 = w_valid_s1_1 & _wen_T_507; // @[Sbuffer.scala 156:25]
  wire  _GEN_12176 = 4'h0 == w_addr_s1_1 | _GEN_8112; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12177 = 4'h1 == w_addr_s1_1 | _GEN_8113; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12178 = 4'h2 == w_addr_s1_1 | _GEN_8114; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12179 = 4'h3 == w_addr_s1_1 | _GEN_8115; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12180 = 4'h4 == w_addr_s1_1 | _GEN_8116; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12181 = 4'h5 == w_addr_s1_1 | _GEN_8117; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12182 = 4'h6 == w_addr_s1_1 | _GEN_8118; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12183 = 4'h7 == w_addr_s1_1 | _GEN_8119; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12184 = 4'h8 == w_addr_s1_1 | _GEN_8120; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12185 = 4'h9 == w_addr_s1_1 | _GEN_8121; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12186 = 4'ha == w_addr_s1_1 | _GEN_8122; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12187 = 4'hb == w_addr_s1_1 | _GEN_8123; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12188 = 4'hc == w_addr_s1_1 | _GEN_8124; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12189 = 4'hd == w_addr_s1_1 | _GEN_8125; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12190 = 4'he == w_addr_s1_1 | _GEN_8126; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12191 = 4'hf == w_addr_s1_1 | _GEN_8127; // @[Sbuffer.scala 162:{42,42}]
  wire  _wen_T_511 = w_mask_s1_1[7] & w_word_offset_s1_1 == 3'h7 | w_wline_s1_1; // @[Sbuffer.scala 157:70]
  wire  wen_127 = w_valid_s1_1 & _wen_T_511; // @[Sbuffer.scala 156:25]
  wire  _GEN_12240 = 4'h0 == w_addr_s1_1 | _GEN_8176; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12241 = 4'h1 == w_addr_s1_1 | _GEN_8177; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12242 = 4'h2 == w_addr_s1_1 | _GEN_8178; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12243 = 4'h3 == w_addr_s1_1 | _GEN_8179; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12244 = 4'h4 == w_addr_s1_1 | _GEN_8180; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12245 = 4'h5 == w_addr_s1_1 | _GEN_8181; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12246 = 4'h6 == w_addr_s1_1 | _GEN_8182; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12247 = 4'h7 == w_addr_s1_1 | _GEN_8183; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12248 = 4'h8 == w_addr_s1_1 | _GEN_8184; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12249 = 4'h9 == w_addr_s1_1 | _GEN_8185; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12250 = 4'ha == w_addr_s1_1 | _GEN_8186; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12251 = 4'hb == w_addr_s1_1 | _GEN_8187; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12252 = 4'hc == w_addr_s1_1 | _GEN_8188; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12253 = 4'hd == w_addr_s1_1 | _GEN_8189; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12254 = 4'he == w_addr_s1_1 | _GEN_8190; // @[Sbuffer.scala 162:{42,42}]
  wire  _GEN_12255 = 4'hf == w_addr_s1_1 | _GEN_8191; // @[Sbuffer.scala 162:{42,42}]
  assign io_dataOut_0_0_0 = data_0_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_1 = data_0_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_2 = data_0_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_3 = data_0_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_4 = data_0_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_5 = data_0_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_6 = data_0_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_0_7 = data_0_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_0 = data_0_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_1 = data_0_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_2 = data_0_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_3 = data_0_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_4 = data_0_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_5 = data_0_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_6 = data_0_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_1_7 = data_0_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_0 = data_0_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_1 = data_0_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_2 = data_0_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_3 = data_0_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_4 = data_0_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_5 = data_0_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_6 = data_0_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_2_7 = data_0_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_0 = data_0_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_1 = data_0_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_2 = data_0_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_3 = data_0_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_4 = data_0_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_5 = data_0_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_6 = data_0_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_3_7 = data_0_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_0 = data_0_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_1 = data_0_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_2 = data_0_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_3 = data_0_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_4 = data_0_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_5 = data_0_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_6 = data_0_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_4_7 = data_0_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_0 = data_0_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_1 = data_0_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_2 = data_0_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_3 = data_0_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_4 = data_0_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_5 = data_0_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_6 = data_0_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_5_7 = data_0_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_0 = data_0_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_1 = data_0_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_2 = data_0_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_3 = data_0_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_4 = data_0_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_5 = data_0_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_6 = data_0_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_6_7 = data_0_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_0 = data_0_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_1 = data_0_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_2 = data_0_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_3 = data_0_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_4 = data_0_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_5 = data_0_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_6 = data_0_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_0_7_7 = data_0_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_0 = data_1_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_1 = data_1_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_2 = data_1_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_3 = data_1_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_4 = data_1_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_5 = data_1_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_6 = data_1_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_0_7 = data_1_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_0 = data_1_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_1 = data_1_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_2 = data_1_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_3 = data_1_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_4 = data_1_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_5 = data_1_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_6 = data_1_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_1_7 = data_1_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_0 = data_1_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_1 = data_1_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_2 = data_1_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_3 = data_1_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_4 = data_1_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_5 = data_1_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_6 = data_1_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_2_7 = data_1_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_0 = data_1_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_1 = data_1_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_2 = data_1_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_3 = data_1_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_4 = data_1_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_5 = data_1_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_6 = data_1_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_3_7 = data_1_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_0 = data_1_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_1 = data_1_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_2 = data_1_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_3 = data_1_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_4 = data_1_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_5 = data_1_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_6 = data_1_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_4_7 = data_1_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_0 = data_1_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_1 = data_1_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_2 = data_1_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_3 = data_1_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_4 = data_1_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_5 = data_1_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_6 = data_1_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_5_7 = data_1_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_0 = data_1_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_1 = data_1_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_2 = data_1_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_3 = data_1_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_4 = data_1_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_5 = data_1_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_6 = data_1_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_6_7 = data_1_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_0 = data_1_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_1 = data_1_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_2 = data_1_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_3 = data_1_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_4 = data_1_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_5 = data_1_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_6 = data_1_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_1_7_7 = data_1_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_0 = data_2_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_1 = data_2_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_2 = data_2_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_3 = data_2_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_4 = data_2_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_5 = data_2_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_6 = data_2_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_0_7 = data_2_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_0 = data_2_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_1 = data_2_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_2 = data_2_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_3 = data_2_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_4 = data_2_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_5 = data_2_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_6 = data_2_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_1_7 = data_2_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_0 = data_2_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_1 = data_2_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_2 = data_2_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_3 = data_2_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_4 = data_2_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_5 = data_2_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_6 = data_2_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_2_7 = data_2_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_0 = data_2_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_1 = data_2_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_2 = data_2_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_3 = data_2_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_4 = data_2_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_5 = data_2_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_6 = data_2_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_3_7 = data_2_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_0 = data_2_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_1 = data_2_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_2 = data_2_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_3 = data_2_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_4 = data_2_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_5 = data_2_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_6 = data_2_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_4_7 = data_2_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_0 = data_2_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_1 = data_2_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_2 = data_2_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_3 = data_2_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_4 = data_2_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_5 = data_2_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_6 = data_2_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_5_7 = data_2_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_0 = data_2_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_1 = data_2_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_2 = data_2_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_3 = data_2_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_4 = data_2_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_5 = data_2_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_6 = data_2_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_6_7 = data_2_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_0 = data_2_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_1 = data_2_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_2 = data_2_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_3 = data_2_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_4 = data_2_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_5 = data_2_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_6 = data_2_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_2_7_7 = data_2_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_0 = data_3_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_1 = data_3_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_2 = data_3_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_3 = data_3_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_4 = data_3_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_5 = data_3_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_6 = data_3_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_0_7 = data_3_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_0 = data_3_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_1 = data_3_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_2 = data_3_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_3 = data_3_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_4 = data_3_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_5 = data_3_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_6 = data_3_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_1_7 = data_3_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_0 = data_3_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_1 = data_3_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_2 = data_3_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_3 = data_3_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_4 = data_3_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_5 = data_3_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_6 = data_3_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_2_7 = data_3_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_0 = data_3_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_1 = data_3_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_2 = data_3_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_3 = data_3_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_4 = data_3_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_5 = data_3_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_6 = data_3_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_3_7 = data_3_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_0 = data_3_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_1 = data_3_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_2 = data_3_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_3 = data_3_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_4 = data_3_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_5 = data_3_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_6 = data_3_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_4_7 = data_3_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_0 = data_3_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_1 = data_3_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_2 = data_3_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_3 = data_3_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_4 = data_3_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_5 = data_3_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_6 = data_3_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_5_7 = data_3_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_0 = data_3_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_1 = data_3_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_2 = data_3_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_3 = data_3_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_4 = data_3_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_5 = data_3_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_6 = data_3_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_6_7 = data_3_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_0 = data_3_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_1 = data_3_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_2 = data_3_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_3 = data_3_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_4 = data_3_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_5 = data_3_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_6 = data_3_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_3_7_7 = data_3_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_0 = data_4_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_1 = data_4_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_2 = data_4_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_3 = data_4_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_4 = data_4_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_5 = data_4_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_6 = data_4_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_0_7 = data_4_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_0 = data_4_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_1 = data_4_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_2 = data_4_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_3 = data_4_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_4 = data_4_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_5 = data_4_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_6 = data_4_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_1_7 = data_4_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_0 = data_4_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_1 = data_4_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_2 = data_4_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_3 = data_4_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_4 = data_4_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_5 = data_4_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_6 = data_4_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_2_7 = data_4_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_0 = data_4_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_1 = data_4_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_2 = data_4_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_3 = data_4_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_4 = data_4_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_5 = data_4_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_6 = data_4_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_3_7 = data_4_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_0 = data_4_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_1 = data_4_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_2 = data_4_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_3 = data_4_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_4 = data_4_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_5 = data_4_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_6 = data_4_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_4_7 = data_4_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_0 = data_4_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_1 = data_4_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_2 = data_4_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_3 = data_4_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_4 = data_4_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_5 = data_4_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_6 = data_4_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_5_7 = data_4_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_0 = data_4_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_1 = data_4_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_2 = data_4_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_3 = data_4_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_4 = data_4_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_5 = data_4_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_6 = data_4_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_6_7 = data_4_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_0 = data_4_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_1 = data_4_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_2 = data_4_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_3 = data_4_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_4 = data_4_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_5 = data_4_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_6 = data_4_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_4_7_7 = data_4_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_0 = data_5_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_1 = data_5_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_2 = data_5_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_3 = data_5_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_4 = data_5_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_5 = data_5_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_6 = data_5_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_0_7 = data_5_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_0 = data_5_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_1 = data_5_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_2 = data_5_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_3 = data_5_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_4 = data_5_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_5 = data_5_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_6 = data_5_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_1_7 = data_5_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_0 = data_5_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_1 = data_5_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_2 = data_5_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_3 = data_5_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_4 = data_5_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_5 = data_5_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_6 = data_5_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_2_7 = data_5_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_0 = data_5_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_1 = data_5_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_2 = data_5_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_3 = data_5_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_4 = data_5_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_5 = data_5_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_6 = data_5_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_3_7 = data_5_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_0 = data_5_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_1 = data_5_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_2 = data_5_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_3 = data_5_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_4 = data_5_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_5 = data_5_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_6 = data_5_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_4_7 = data_5_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_0 = data_5_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_1 = data_5_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_2 = data_5_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_3 = data_5_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_4 = data_5_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_5 = data_5_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_6 = data_5_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_5_7 = data_5_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_0 = data_5_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_1 = data_5_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_2 = data_5_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_3 = data_5_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_4 = data_5_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_5 = data_5_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_6 = data_5_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_6_7 = data_5_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_0 = data_5_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_1 = data_5_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_2 = data_5_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_3 = data_5_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_4 = data_5_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_5 = data_5_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_6 = data_5_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_5_7_7 = data_5_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_0 = data_6_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_1 = data_6_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_2 = data_6_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_3 = data_6_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_4 = data_6_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_5 = data_6_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_6 = data_6_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_0_7 = data_6_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_0 = data_6_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_1 = data_6_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_2 = data_6_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_3 = data_6_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_4 = data_6_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_5 = data_6_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_6 = data_6_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_1_7 = data_6_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_0 = data_6_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_1 = data_6_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_2 = data_6_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_3 = data_6_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_4 = data_6_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_5 = data_6_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_6 = data_6_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_2_7 = data_6_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_0 = data_6_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_1 = data_6_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_2 = data_6_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_3 = data_6_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_4 = data_6_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_5 = data_6_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_6 = data_6_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_3_7 = data_6_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_0 = data_6_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_1 = data_6_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_2 = data_6_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_3 = data_6_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_4 = data_6_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_5 = data_6_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_6 = data_6_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_4_7 = data_6_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_0 = data_6_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_1 = data_6_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_2 = data_6_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_3 = data_6_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_4 = data_6_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_5 = data_6_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_6 = data_6_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_5_7 = data_6_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_0 = data_6_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_1 = data_6_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_2 = data_6_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_3 = data_6_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_4 = data_6_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_5 = data_6_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_6 = data_6_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_6_7 = data_6_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_0 = data_6_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_1 = data_6_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_2 = data_6_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_3 = data_6_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_4 = data_6_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_5 = data_6_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_6 = data_6_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_6_7_7 = data_6_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_0 = data_7_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_1 = data_7_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_2 = data_7_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_3 = data_7_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_4 = data_7_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_5 = data_7_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_6 = data_7_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_0_7 = data_7_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_0 = data_7_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_1 = data_7_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_2 = data_7_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_3 = data_7_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_4 = data_7_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_5 = data_7_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_6 = data_7_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_1_7 = data_7_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_0 = data_7_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_1 = data_7_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_2 = data_7_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_3 = data_7_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_4 = data_7_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_5 = data_7_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_6 = data_7_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_2_7 = data_7_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_0 = data_7_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_1 = data_7_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_2 = data_7_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_3 = data_7_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_4 = data_7_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_5 = data_7_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_6 = data_7_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_3_7 = data_7_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_0 = data_7_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_1 = data_7_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_2 = data_7_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_3 = data_7_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_4 = data_7_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_5 = data_7_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_6 = data_7_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_4_7 = data_7_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_0 = data_7_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_1 = data_7_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_2 = data_7_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_3 = data_7_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_4 = data_7_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_5 = data_7_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_6 = data_7_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_5_7 = data_7_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_0 = data_7_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_1 = data_7_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_2 = data_7_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_3 = data_7_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_4 = data_7_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_5 = data_7_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_6 = data_7_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_6_7 = data_7_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_0 = data_7_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_1 = data_7_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_2 = data_7_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_3 = data_7_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_4 = data_7_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_5 = data_7_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_6 = data_7_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_7_7_7 = data_7_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_0 = data_8_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_1 = data_8_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_2 = data_8_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_3 = data_8_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_4 = data_8_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_5 = data_8_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_6 = data_8_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_0_7 = data_8_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_0 = data_8_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_1 = data_8_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_2 = data_8_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_3 = data_8_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_4 = data_8_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_5 = data_8_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_6 = data_8_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_1_7 = data_8_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_0 = data_8_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_1 = data_8_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_2 = data_8_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_3 = data_8_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_4 = data_8_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_5 = data_8_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_6 = data_8_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_2_7 = data_8_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_0 = data_8_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_1 = data_8_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_2 = data_8_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_3 = data_8_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_4 = data_8_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_5 = data_8_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_6 = data_8_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_3_7 = data_8_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_0 = data_8_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_1 = data_8_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_2 = data_8_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_3 = data_8_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_4 = data_8_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_5 = data_8_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_6 = data_8_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_4_7 = data_8_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_0 = data_8_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_1 = data_8_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_2 = data_8_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_3 = data_8_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_4 = data_8_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_5 = data_8_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_6 = data_8_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_5_7 = data_8_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_0 = data_8_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_1 = data_8_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_2 = data_8_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_3 = data_8_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_4 = data_8_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_5 = data_8_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_6 = data_8_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_6_7 = data_8_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_0 = data_8_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_1 = data_8_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_2 = data_8_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_3 = data_8_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_4 = data_8_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_5 = data_8_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_6 = data_8_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_8_7_7 = data_8_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_0 = data_9_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_1 = data_9_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_2 = data_9_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_3 = data_9_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_4 = data_9_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_5 = data_9_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_6 = data_9_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_0_7 = data_9_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_0 = data_9_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_1 = data_9_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_2 = data_9_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_3 = data_9_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_4 = data_9_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_5 = data_9_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_6 = data_9_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_1_7 = data_9_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_0 = data_9_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_1 = data_9_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_2 = data_9_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_3 = data_9_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_4 = data_9_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_5 = data_9_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_6 = data_9_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_2_7 = data_9_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_0 = data_9_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_1 = data_9_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_2 = data_9_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_3 = data_9_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_4 = data_9_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_5 = data_9_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_6 = data_9_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_3_7 = data_9_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_0 = data_9_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_1 = data_9_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_2 = data_9_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_3 = data_9_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_4 = data_9_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_5 = data_9_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_6 = data_9_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_4_7 = data_9_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_0 = data_9_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_1 = data_9_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_2 = data_9_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_3 = data_9_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_4 = data_9_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_5 = data_9_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_6 = data_9_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_5_7 = data_9_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_0 = data_9_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_1 = data_9_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_2 = data_9_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_3 = data_9_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_4 = data_9_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_5 = data_9_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_6 = data_9_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_6_7 = data_9_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_0 = data_9_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_1 = data_9_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_2 = data_9_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_3 = data_9_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_4 = data_9_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_5 = data_9_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_6 = data_9_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_9_7_7 = data_9_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_0 = data_10_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_1 = data_10_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_2 = data_10_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_3 = data_10_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_4 = data_10_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_5 = data_10_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_6 = data_10_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_0_7 = data_10_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_0 = data_10_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_1 = data_10_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_2 = data_10_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_3 = data_10_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_4 = data_10_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_5 = data_10_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_6 = data_10_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_1_7 = data_10_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_0 = data_10_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_1 = data_10_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_2 = data_10_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_3 = data_10_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_4 = data_10_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_5 = data_10_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_6 = data_10_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_2_7 = data_10_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_0 = data_10_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_1 = data_10_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_2 = data_10_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_3 = data_10_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_4 = data_10_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_5 = data_10_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_6 = data_10_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_3_7 = data_10_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_0 = data_10_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_1 = data_10_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_2 = data_10_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_3 = data_10_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_4 = data_10_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_5 = data_10_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_6 = data_10_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_4_7 = data_10_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_0 = data_10_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_1 = data_10_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_2 = data_10_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_3 = data_10_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_4 = data_10_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_5 = data_10_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_6 = data_10_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_5_7 = data_10_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_0 = data_10_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_1 = data_10_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_2 = data_10_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_3 = data_10_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_4 = data_10_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_5 = data_10_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_6 = data_10_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_6_7 = data_10_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_0 = data_10_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_1 = data_10_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_2 = data_10_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_3 = data_10_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_4 = data_10_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_5 = data_10_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_6 = data_10_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_10_7_7 = data_10_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_0 = data_11_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_1 = data_11_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_2 = data_11_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_3 = data_11_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_4 = data_11_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_5 = data_11_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_6 = data_11_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_0_7 = data_11_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_0 = data_11_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_1 = data_11_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_2 = data_11_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_3 = data_11_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_4 = data_11_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_5 = data_11_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_6 = data_11_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_1_7 = data_11_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_0 = data_11_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_1 = data_11_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_2 = data_11_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_3 = data_11_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_4 = data_11_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_5 = data_11_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_6 = data_11_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_2_7 = data_11_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_0 = data_11_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_1 = data_11_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_2 = data_11_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_3 = data_11_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_4 = data_11_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_5 = data_11_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_6 = data_11_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_3_7 = data_11_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_0 = data_11_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_1 = data_11_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_2 = data_11_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_3 = data_11_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_4 = data_11_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_5 = data_11_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_6 = data_11_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_4_7 = data_11_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_0 = data_11_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_1 = data_11_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_2 = data_11_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_3 = data_11_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_4 = data_11_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_5 = data_11_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_6 = data_11_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_5_7 = data_11_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_0 = data_11_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_1 = data_11_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_2 = data_11_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_3 = data_11_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_4 = data_11_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_5 = data_11_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_6 = data_11_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_6_7 = data_11_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_0 = data_11_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_1 = data_11_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_2 = data_11_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_3 = data_11_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_4 = data_11_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_5 = data_11_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_6 = data_11_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_11_7_7 = data_11_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_0 = data_12_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_1 = data_12_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_2 = data_12_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_3 = data_12_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_4 = data_12_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_5 = data_12_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_6 = data_12_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_0_7 = data_12_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_0 = data_12_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_1 = data_12_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_2 = data_12_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_3 = data_12_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_4 = data_12_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_5 = data_12_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_6 = data_12_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_1_7 = data_12_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_0 = data_12_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_1 = data_12_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_2 = data_12_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_3 = data_12_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_4 = data_12_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_5 = data_12_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_6 = data_12_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_2_7 = data_12_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_0 = data_12_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_1 = data_12_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_2 = data_12_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_3 = data_12_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_4 = data_12_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_5 = data_12_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_6 = data_12_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_3_7 = data_12_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_0 = data_12_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_1 = data_12_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_2 = data_12_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_3 = data_12_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_4 = data_12_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_5 = data_12_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_6 = data_12_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_4_7 = data_12_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_0 = data_12_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_1 = data_12_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_2 = data_12_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_3 = data_12_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_4 = data_12_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_5 = data_12_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_6 = data_12_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_5_7 = data_12_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_0 = data_12_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_1 = data_12_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_2 = data_12_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_3 = data_12_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_4 = data_12_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_5 = data_12_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_6 = data_12_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_6_7 = data_12_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_0 = data_12_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_1 = data_12_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_2 = data_12_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_3 = data_12_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_4 = data_12_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_5 = data_12_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_6 = data_12_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_12_7_7 = data_12_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_0 = data_13_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_1 = data_13_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_2 = data_13_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_3 = data_13_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_4 = data_13_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_5 = data_13_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_6 = data_13_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_0_7 = data_13_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_0 = data_13_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_1 = data_13_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_2 = data_13_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_3 = data_13_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_4 = data_13_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_5 = data_13_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_6 = data_13_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_1_7 = data_13_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_0 = data_13_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_1 = data_13_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_2 = data_13_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_3 = data_13_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_4 = data_13_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_5 = data_13_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_6 = data_13_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_2_7 = data_13_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_0 = data_13_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_1 = data_13_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_2 = data_13_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_3 = data_13_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_4 = data_13_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_5 = data_13_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_6 = data_13_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_3_7 = data_13_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_0 = data_13_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_1 = data_13_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_2 = data_13_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_3 = data_13_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_4 = data_13_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_5 = data_13_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_6 = data_13_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_4_7 = data_13_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_0 = data_13_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_1 = data_13_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_2 = data_13_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_3 = data_13_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_4 = data_13_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_5 = data_13_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_6 = data_13_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_5_7 = data_13_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_0 = data_13_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_1 = data_13_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_2 = data_13_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_3 = data_13_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_4 = data_13_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_5 = data_13_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_6 = data_13_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_6_7 = data_13_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_0 = data_13_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_1 = data_13_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_2 = data_13_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_3 = data_13_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_4 = data_13_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_5 = data_13_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_6 = data_13_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_13_7_7 = data_13_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_0 = data_14_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_1 = data_14_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_2 = data_14_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_3 = data_14_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_4 = data_14_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_5 = data_14_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_6 = data_14_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_0_7 = data_14_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_0 = data_14_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_1 = data_14_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_2 = data_14_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_3 = data_14_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_4 = data_14_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_5 = data_14_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_6 = data_14_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_1_7 = data_14_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_0 = data_14_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_1 = data_14_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_2 = data_14_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_3 = data_14_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_4 = data_14_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_5 = data_14_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_6 = data_14_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_2_7 = data_14_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_0 = data_14_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_1 = data_14_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_2 = data_14_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_3 = data_14_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_4 = data_14_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_5 = data_14_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_6 = data_14_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_3_7 = data_14_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_0 = data_14_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_1 = data_14_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_2 = data_14_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_3 = data_14_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_4 = data_14_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_5 = data_14_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_6 = data_14_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_4_7 = data_14_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_0 = data_14_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_1 = data_14_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_2 = data_14_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_3 = data_14_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_4 = data_14_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_5 = data_14_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_6 = data_14_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_5_7 = data_14_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_0 = data_14_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_1 = data_14_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_2 = data_14_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_3 = data_14_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_4 = data_14_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_5 = data_14_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_6 = data_14_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_6_7 = data_14_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_0 = data_14_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_1 = data_14_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_2 = data_14_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_3 = data_14_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_4 = data_14_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_5 = data_14_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_6 = data_14_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_14_7_7 = data_14_7_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_0 = data_15_0_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_1 = data_15_0_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_2 = data_15_0_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_3 = data_15_0_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_4 = data_15_0_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_5 = data_15_0_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_6 = data_15_0_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_0_7 = data_15_0_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_0 = data_15_1_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_1 = data_15_1_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_2 = data_15_1_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_3 = data_15_1_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_4 = data_15_1_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_5 = data_15_1_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_6 = data_15_1_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_1_7 = data_15_1_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_0 = data_15_2_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_1 = data_15_2_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_2 = data_15_2_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_3 = data_15_2_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_4 = data_15_2_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_5 = data_15_2_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_6 = data_15_2_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_2_7 = data_15_2_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_0 = data_15_3_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_1 = data_15_3_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_2 = data_15_3_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_3 = data_15_3_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_4 = data_15_3_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_5 = data_15_3_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_6 = data_15_3_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_3_7 = data_15_3_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_0 = data_15_4_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_1 = data_15_4_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_2 = data_15_4_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_3 = data_15_4_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_4 = data_15_4_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_5 = data_15_4_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_6 = data_15_4_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_4_7 = data_15_4_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_0 = data_15_5_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_1 = data_15_5_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_2 = data_15_5_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_3 = data_15_5_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_4 = data_15_5_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_5 = data_15_5_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_6 = data_15_5_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_5_7 = data_15_5_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_0 = data_15_6_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_1 = data_15_6_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_2 = data_15_6_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_3 = data_15_6_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_4 = data_15_6_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_5 = data_15_6_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_6 = data_15_6_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_6_7 = data_15_6_7; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_0 = data_15_7_0; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_1 = data_15_7_1; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_2 = data_15_7_2; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_3 = data_15_7_3; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_4 = data_15_7_4; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_5 = data_15_7_5; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_6 = data_15_7_6; // @[Sbuffer.scala 224:14]
  assign io_dataOut_15_7_7 = data_15_7_7; // @[Sbuffer.scala 224:14]
  assign io_maskOut_0_0_0 = mask_0_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_1 = mask_0_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_2 = mask_0_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_3 = mask_0_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_4 = mask_0_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_5 = mask_0_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_6 = mask_0_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_0_7 = mask_0_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_0 = mask_0_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_1 = mask_0_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_2 = mask_0_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_3 = mask_0_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_4 = mask_0_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_5 = mask_0_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_6 = mask_0_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_1_7 = mask_0_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_0 = mask_0_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_1 = mask_0_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_2 = mask_0_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_3 = mask_0_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_4 = mask_0_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_5 = mask_0_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_6 = mask_0_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_2_7 = mask_0_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_0 = mask_0_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_1 = mask_0_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_2 = mask_0_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_3 = mask_0_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_4 = mask_0_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_5 = mask_0_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_6 = mask_0_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_3_7 = mask_0_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_0 = mask_0_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_1 = mask_0_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_2 = mask_0_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_3 = mask_0_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_4 = mask_0_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_5 = mask_0_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_6 = mask_0_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_4_7 = mask_0_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_0 = mask_0_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_1 = mask_0_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_2 = mask_0_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_3 = mask_0_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_4 = mask_0_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_5 = mask_0_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_6 = mask_0_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_5_7 = mask_0_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_0 = mask_0_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_1 = mask_0_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_2 = mask_0_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_3 = mask_0_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_4 = mask_0_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_5 = mask_0_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_6 = mask_0_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_6_7 = mask_0_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_0 = mask_0_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_1 = mask_0_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_2 = mask_0_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_3 = mask_0_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_4 = mask_0_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_5 = mask_0_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_6 = mask_0_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_0_7_7 = mask_0_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_0 = mask_1_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_1 = mask_1_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_2 = mask_1_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_3 = mask_1_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_4 = mask_1_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_5 = mask_1_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_6 = mask_1_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_0_7 = mask_1_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_0 = mask_1_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_1 = mask_1_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_2 = mask_1_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_3 = mask_1_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_4 = mask_1_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_5 = mask_1_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_6 = mask_1_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_1_7 = mask_1_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_0 = mask_1_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_1 = mask_1_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_2 = mask_1_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_3 = mask_1_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_4 = mask_1_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_5 = mask_1_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_6 = mask_1_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_2_7 = mask_1_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_0 = mask_1_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_1 = mask_1_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_2 = mask_1_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_3 = mask_1_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_4 = mask_1_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_5 = mask_1_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_6 = mask_1_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_3_7 = mask_1_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_0 = mask_1_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_1 = mask_1_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_2 = mask_1_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_3 = mask_1_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_4 = mask_1_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_5 = mask_1_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_6 = mask_1_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_4_7 = mask_1_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_0 = mask_1_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_1 = mask_1_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_2 = mask_1_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_3 = mask_1_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_4 = mask_1_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_5 = mask_1_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_6 = mask_1_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_5_7 = mask_1_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_0 = mask_1_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_1 = mask_1_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_2 = mask_1_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_3 = mask_1_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_4 = mask_1_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_5 = mask_1_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_6 = mask_1_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_6_7 = mask_1_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_0 = mask_1_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_1 = mask_1_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_2 = mask_1_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_3 = mask_1_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_4 = mask_1_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_5 = mask_1_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_6 = mask_1_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_1_7_7 = mask_1_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_0 = mask_2_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_1 = mask_2_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_2 = mask_2_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_3 = mask_2_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_4 = mask_2_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_5 = mask_2_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_6 = mask_2_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_0_7 = mask_2_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_0 = mask_2_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_1 = mask_2_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_2 = mask_2_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_3 = mask_2_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_4 = mask_2_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_5 = mask_2_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_6 = mask_2_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_1_7 = mask_2_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_0 = mask_2_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_1 = mask_2_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_2 = mask_2_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_3 = mask_2_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_4 = mask_2_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_5 = mask_2_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_6 = mask_2_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_2_7 = mask_2_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_0 = mask_2_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_1 = mask_2_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_2 = mask_2_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_3 = mask_2_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_4 = mask_2_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_5 = mask_2_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_6 = mask_2_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_3_7 = mask_2_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_0 = mask_2_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_1 = mask_2_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_2 = mask_2_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_3 = mask_2_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_4 = mask_2_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_5 = mask_2_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_6 = mask_2_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_4_7 = mask_2_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_0 = mask_2_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_1 = mask_2_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_2 = mask_2_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_3 = mask_2_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_4 = mask_2_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_5 = mask_2_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_6 = mask_2_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_5_7 = mask_2_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_0 = mask_2_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_1 = mask_2_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_2 = mask_2_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_3 = mask_2_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_4 = mask_2_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_5 = mask_2_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_6 = mask_2_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_6_7 = mask_2_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_0 = mask_2_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_1 = mask_2_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_2 = mask_2_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_3 = mask_2_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_4 = mask_2_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_5 = mask_2_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_6 = mask_2_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_2_7_7 = mask_2_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_0 = mask_3_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_1 = mask_3_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_2 = mask_3_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_3 = mask_3_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_4 = mask_3_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_5 = mask_3_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_6 = mask_3_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_0_7 = mask_3_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_0 = mask_3_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_1 = mask_3_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_2 = mask_3_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_3 = mask_3_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_4 = mask_3_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_5 = mask_3_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_6 = mask_3_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_1_7 = mask_3_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_0 = mask_3_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_1 = mask_3_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_2 = mask_3_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_3 = mask_3_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_4 = mask_3_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_5 = mask_3_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_6 = mask_3_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_2_7 = mask_3_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_0 = mask_3_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_1 = mask_3_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_2 = mask_3_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_3 = mask_3_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_4 = mask_3_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_5 = mask_3_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_6 = mask_3_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_3_7 = mask_3_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_0 = mask_3_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_1 = mask_3_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_2 = mask_3_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_3 = mask_3_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_4 = mask_3_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_5 = mask_3_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_6 = mask_3_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_4_7 = mask_3_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_0 = mask_3_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_1 = mask_3_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_2 = mask_3_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_3 = mask_3_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_4 = mask_3_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_5 = mask_3_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_6 = mask_3_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_5_7 = mask_3_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_0 = mask_3_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_1 = mask_3_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_2 = mask_3_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_3 = mask_3_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_4 = mask_3_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_5 = mask_3_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_6 = mask_3_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_6_7 = mask_3_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_0 = mask_3_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_1 = mask_3_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_2 = mask_3_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_3 = mask_3_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_4 = mask_3_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_5 = mask_3_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_6 = mask_3_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_3_7_7 = mask_3_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_0 = mask_4_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_1 = mask_4_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_2 = mask_4_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_3 = mask_4_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_4 = mask_4_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_5 = mask_4_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_6 = mask_4_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_0_7 = mask_4_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_0 = mask_4_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_1 = mask_4_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_2 = mask_4_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_3 = mask_4_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_4 = mask_4_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_5 = mask_4_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_6 = mask_4_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_1_7 = mask_4_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_0 = mask_4_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_1 = mask_4_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_2 = mask_4_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_3 = mask_4_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_4 = mask_4_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_5 = mask_4_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_6 = mask_4_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_2_7 = mask_4_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_0 = mask_4_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_1 = mask_4_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_2 = mask_4_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_3 = mask_4_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_4 = mask_4_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_5 = mask_4_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_6 = mask_4_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_3_7 = mask_4_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_0 = mask_4_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_1 = mask_4_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_2 = mask_4_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_3 = mask_4_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_4 = mask_4_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_5 = mask_4_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_6 = mask_4_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_4_7 = mask_4_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_0 = mask_4_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_1 = mask_4_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_2 = mask_4_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_3 = mask_4_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_4 = mask_4_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_5 = mask_4_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_6 = mask_4_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_5_7 = mask_4_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_0 = mask_4_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_1 = mask_4_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_2 = mask_4_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_3 = mask_4_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_4 = mask_4_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_5 = mask_4_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_6 = mask_4_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_6_7 = mask_4_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_0 = mask_4_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_1 = mask_4_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_2 = mask_4_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_3 = mask_4_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_4 = mask_4_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_5 = mask_4_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_6 = mask_4_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_4_7_7 = mask_4_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_0 = mask_5_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_1 = mask_5_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_2 = mask_5_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_3 = mask_5_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_4 = mask_5_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_5 = mask_5_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_6 = mask_5_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_0_7 = mask_5_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_0 = mask_5_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_1 = mask_5_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_2 = mask_5_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_3 = mask_5_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_4 = mask_5_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_5 = mask_5_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_6 = mask_5_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_1_7 = mask_5_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_0 = mask_5_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_1 = mask_5_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_2 = mask_5_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_3 = mask_5_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_4 = mask_5_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_5 = mask_5_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_6 = mask_5_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_2_7 = mask_5_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_0 = mask_5_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_1 = mask_5_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_2 = mask_5_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_3 = mask_5_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_4 = mask_5_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_5 = mask_5_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_6 = mask_5_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_3_7 = mask_5_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_0 = mask_5_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_1 = mask_5_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_2 = mask_5_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_3 = mask_5_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_4 = mask_5_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_5 = mask_5_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_6 = mask_5_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_4_7 = mask_5_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_0 = mask_5_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_1 = mask_5_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_2 = mask_5_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_3 = mask_5_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_4 = mask_5_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_5 = mask_5_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_6 = mask_5_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_5_7 = mask_5_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_0 = mask_5_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_1 = mask_5_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_2 = mask_5_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_3 = mask_5_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_4 = mask_5_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_5 = mask_5_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_6 = mask_5_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_6_7 = mask_5_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_0 = mask_5_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_1 = mask_5_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_2 = mask_5_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_3 = mask_5_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_4 = mask_5_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_5 = mask_5_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_6 = mask_5_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_5_7_7 = mask_5_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_0 = mask_6_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_1 = mask_6_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_2 = mask_6_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_3 = mask_6_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_4 = mask_6_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_5 = mask_6_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_6 = mask_6_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_0_7 = mask_6_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_0 = mask_6_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_1 = mask_6_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_2 = mask_6_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_3 = mask_6_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_4 = mask_6_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_5 = mask_6_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_6 = mask_6_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_1_7 = mask_6_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_0 = mask_6_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_1 = mask_6_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_2 = mask_6_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_3 = mask_6_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_4 = mask_6_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_5 = mask_6_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_6 = mask_6_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_2_7 = mask_6_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_0 = mask_6_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_1 = mask_6_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_2 = mask_6_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_3 = mask_6_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_4 = mask_6_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_5 = mask_6_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_6 = mask_6_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_3_7 = mask_6_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_0 = mask_6_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_1 = mask_6_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_2 = mask_6_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_3 = mask_6_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_4 = mask_6_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_5 = mask_6_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_6 = mask_6_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_4_7 = mask_6_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_0 = mask_6_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_1 = mask_6_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_2 = mask_6_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_3 = mask_6_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_4 = mask_6_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_5 = mask_6_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_6 = mask_6_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_5_7 = mask_6_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_0 = mask_6_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_1 = mask_6_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_2 = mask_6_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_3 = mask_6_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_4 = mask_6_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_5 = mask_6_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_6 = mask_6_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_6_7 = mask_6_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_0 = mask_6_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_1 = mask_6_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_2 = mask_6_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_3 = mask_6_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_4 = mask_6_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_5 = mask_6_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_6 = mask_6_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_6_7_7 = mask_6_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_0 = mask_7_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_1 = mask_7_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_2 = mask_7_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_3 = mask_7_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_4 = mask_7_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_5 = mask_7_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_6 = mask_7_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_0_7 = mask_7_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_0 = mask_7_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_1 = mask_7_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_2 = mask_7_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_3 = mask_7_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_4 = mask_7_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_5 = mask_7_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_6 = mask_7_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_1_7 = mask_7_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_0 = mask_7_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_1 = mask_7_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_2 = mask_7_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_3 = mask_7_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_4 = mask_7_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_5 = mask_7_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_6 = mask_7_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_2_7 = mask_7_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_0 = mask_7_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_1 = mask_7_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_2 = mask_7_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_3 = mask_7_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_4 = mask_7_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_5 = mask_7_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_6 = mask_7_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_3_7 = mask_7_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_0 = mask_7_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_1 = mask_7_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_2 = mask_7_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_3 = mask_7_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_4 = mask_7_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_5 = mask_7_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_6 = mask_7_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_4_7 = mask_7_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_0 = mask_7_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_1 = mask_7_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_2 = mask_7_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_3 = mask_7_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_4 = mask_7_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_5 = mask_7_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_6 = mask_7_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_5_7 = mask_7_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_0 = mask_7_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_1 = mask_7_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_2 = mask_7_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_3 = mask_7_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_4 = mask_7_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_5 = mask_7_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_6 = mask_7_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_6_7 = mask_7_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_0 = mask_7_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_1 = mask_7_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_2 = mask_7_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_3 = mask_7_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_4 = mask_7_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_5 = mask_7_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_6 = mask_7_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_7_7_7 = mask_7_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_0 = mask_8_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_1 = mask_8_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_2 = mask_8_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_3 = mask_8_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_4 = mask_8_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_5 = mask_8_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_6 = mask_8_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_0_7 = mask_8_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_0 = mask_8_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_1 = mask_8_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_2 = mask_8_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_3 = mask_8_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_4 = mask_8_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_5 = mask_8_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_6 = mask_8_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_1_7 = mask_8_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_0 = mask_8_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_1 = mask_8_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_2 = mask_8_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_3 = mask_8_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_4 = mask_8_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_5 = mask_8_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_6 = mask_8_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_2_7 = mask_8_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_0 = mask_8_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_1 = mask_8_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_2 = mask_8_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_3 = mask_8_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_4 = mask_8_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_5 = mask_8_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_6 = mask_8_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_3_7 = mask_8_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_0 = mask_8_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_1 = mask_8_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_2 = mask_8_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_3 = mask_8_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_4 = mask_8_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_5 = mask_8_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_6 = mask_8_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_4_7 = mask_8_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_0 = mask_8_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_1 = mask_8_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_2 = mask_8_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_3 = mask_8_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_4 = mask_8_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_5 = mask_8_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_6 = mask_8_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_5_7 = mask_8_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_0 = mask_8_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_1 = mask_8_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_2 = mask_8_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_3 = mask_8_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_4 = mask_8_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_5 = mask_8_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_6 = mask_8_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_6_7 = mask_8_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_0 = mask_8_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_1 = mask_8_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_2 = mask_8_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_3 = mask_8_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_4 = mask_8_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_5 = mask_8_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_6 = mask_8_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_8_7_7 = mask_8_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_0 = mask_9_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_1 = mask_9_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_2 = mask_9_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_3 = mask_9_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_4 = mask_9_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_5 = mask_9_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_6 = mask_9_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_0_7 = mask_9_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_0 = mask_9_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_1 = mask_9_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_2 = mask_9_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_3 = mask_9_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_4 = mask_9_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_5 = mask_9_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_6 = mask_9_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_1_7 = mask_9_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_0 = mask_9_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_1 = mask_9_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_2 = mask_9_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_3 = mask_9_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_4 = mask_9_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_5 = mask_9_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_6 = mask_9_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_2_7 = mask_9_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_0 = mask_9_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_1 = mask_9_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_2 = mask_9_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_3 = mask_9_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_4 = mask_9_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_5 = mask_9_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_6 = mask_9_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_3_7 = mask_9_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_0 = mask_9_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_1 = mask_9_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_2 = mask_9_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_3 = mask_9_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_4 = mask_9_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_5 = mask_9_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_6 = mask_9_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_4_7 = mask_9_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_0 = mask_9_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_1 = mask_9_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_2 = mask_9_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_3 = mask_9_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_4 = mask_9_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_5 = mask_9_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_6 = mask_9_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_5_7 = mask_9_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_0 = mask_9_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_1 = mask_9_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_2 = mask_9_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_3 = mask_9_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_4 = mask_9_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_5 = mask_9_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_6 = mask_9_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_6_7 = mask_9_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_0 = mask_9_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_1 = mask_9_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_2 = mask_9_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_3 = mask_9_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_4 = mask_9_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_5 = mask_9_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_6 = mask_9_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_9_7_7 = mask_9_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_0 = mask_10_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_1 = mask_10_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_2 = mask_10_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_3 = mask_10_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_4 = mask_10_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_5 = mask_10_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_6 = mask_10_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_0_7 = mask_10_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_0 = mask_10_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_1 = mask_10_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_2 = mask_10_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_3 = mask_10_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_4 = mask_10_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_5 = mask_10_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_6 = mask_10_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_1_7 = mask_10_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_0 = mask_10_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_1 = mask_10_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_2 = mask_10_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_3 = mask_10_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_4 = mask_10_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_5 = mask_10_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_6 = mask_10_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_2_7 = mask_10_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_0 = mask_10_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_1 = mask_10_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_2 = mask_10_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_3 = mask_10_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_4 = mask_10_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_5 = mask_10_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_6 = mask_10_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_3_7 = mask_10_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_0 = mask_10_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_1 = mask_10_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_2 = mask_10_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_3 = mask_10_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_4 = mask_10_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_5 = mask_10_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_6 = mask_10_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_4_7 = mask_10_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_0 = mask_10_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_1 = mask_10_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_2 = mask_10_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_3 = mask_10_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_4 = mask_10_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_5 = mask_10_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_6 = mask_10_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_5_7 = mask_10_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_0 = mask_10_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_1 = mask_10_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_2 = mask_10_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_3 = mask_10_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_4 = mask_10_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_5 = mask_10_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_6 = mask_10_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_6_7 = mask_10_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_0 = mask_10_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_1 = mask_10_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_2 = mask_10_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_3 = mask_10_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_4 = mask_10_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_5 = mask_10_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_6 = mask_10_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_10_7_7 = mask_10_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_0 = mask_11_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_1 = mask_11_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_2 = mask_11_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_3 = mask_11_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_4 = mask_11_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_5 = mask_11_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_6 = mask_11_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_0_7 = mask_11_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_0 = mask_11_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_1 = mask_11_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_2 = mask_11_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_3 = mask_11_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_4 = mask_11_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_5 = mask_11_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_6 = mask_11_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_1_7 = mask_11_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_0 = mask_11_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_1 = mask_11_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_2 = mask_11_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_3 = mask_11_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_4 = mask_11_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_5 = mask_11_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_6 = mask_11_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_2_7 = mask_11_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_0 = mask_11_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_1 = mask_11_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_2 = mask_11_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_3 = mask_11_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_4 = mask_11_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_5 = mask_11_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_6 = mask_11_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_3_7 = mask_11_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_0 = mask_11_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_1 = mask_11_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_2 = mask_11_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_3 = mask_11_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_4 = mask_11_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_5 = mask_11_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_6 = mask_11_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_4_7 = mask_11_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_0 = mask_11_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_1 = mask_11_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_2 = mask_11_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_3 = mask_11_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_4 = mask_11_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_5 = mask_11_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_6 = mask_11_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_5_7 = mask_11_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_0 = mask_11_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_1 = mask_11_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_2 = mask_11_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_3 = mask_11_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_4 = mask_11_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_5 = mask_11_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_6 = mask_11_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_6_7 = mask_11_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_0 = mask_11_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_1 = mask_11_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_2 = mask_11_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_3 = mask_11_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_4 = mask_11_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_5 = mask_11_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_6 = mask_11_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_11_7_7 = mask_11_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_0 = mask_12_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_1 = mask_12_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_2 = mask_12_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_3 = mask_12_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_4 = mask_12_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_5 = mask_12_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_6 = mask_12_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_0_7 = mask_12_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_0 = mask_12_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_1 = mask_12_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_2 = mask_12_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_3 = mask_12_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_4 = mask_12_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_5 = mask_12_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_6 = mask_12_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_1_7 = mask_12_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_0 = mask_12_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_1 = mask_12_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_2 = mask_12_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_3 = mask_12_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_4 = mask_12_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_5 = mask_12_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_6 = mask_12_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_2_7 = mask_12_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_0 = mask_12_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_1 = mask_12_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_2 = mask_12_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_3 = mask_12_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_4 = mask_12_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_5 = mask_12_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_6 = mask_12_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_3_7 = mask_12_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_0 = mask_12_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_1 = mask_12_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_2 = mask_12_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_3 = mask_12_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_4 = mask_12_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_5 = mask_12_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_6 = mask_12_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_4_7 = mask_12_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_0 = mask_12_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_1 = mask_12_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_2 = mask_12_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_3 = mask_12_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_4 = mask_12_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_5 = mask_12_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_6 = mask_12_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_5_7 = mask_12_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_0 = mask_12_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_1 = mask_12_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_2 = mask_12_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_3 = mask_12_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_4 = mask_12_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_5 = mask_12_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_6 = mask_12_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_6_7 = mask_12_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_0 = mask_12_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_1 = mask_12_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_2 = mask_12_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_3 = mask_12_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_4 = mask_12_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_5 = mask_12_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_6 = mask_12_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_12_7_7 = mask_12_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_0 = mask_13_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_1 = mask_13_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_2 = mask_13_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_3 = mask_13_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_4 = mask_13_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_5 = mask_13_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_6 = mask_13_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_0_7 = mask_13_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_0 = mask_13_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_1 = mask_13_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_2 = mask_13_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_3 = mask_13_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_4 = mask_13_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_5 = mask_13_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_6 = mask_13_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_1_7 = mask_13_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_0 = mask_13_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_1 = mask_13_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_2 = mask_13_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_3 = mask_13_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_4 = mask_13_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_5 = mask_13_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_6 = mask_13_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_2_7 = mask_13_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_0 = mask_13_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_1 = mask_13_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_2 = mask_13_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_3 = mask_13_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_4 = mask_13_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_5 = mask_13_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_6 = mask_13_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_3_7 = mask_13_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_0 = mask_13_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_1 = mask_13_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_2 = mask_13_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_3 = mask_13_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_4 = mask_13_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_5 = mask_13_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_6 = mask_13_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_4_7 = mask_13_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_0 = mask_13_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_1 = mask_13_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_2 = mask_13_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_3 = mask_13_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_4 = mask_13_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_5 = mask_13_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_6 = mask_13_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_5_7 = mask_13_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_0 = mask_13_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_1 = mask_13_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_2 = mask_13_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_3 = mask_13_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_4 = mask_13_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_5 = mask_13_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_6 = mask_13_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_6_7 = mask_13_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_0 = mask_13_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_1 = mask_13_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_2 = mask_13_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_3 = mask_13_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_4 = mask_13_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_5 = mask_13_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_6 = mask_13_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_13_7_7 = mask_13_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_0 = mask_14_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_1 = mask_14_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_2 = mask_14_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_3 = mask_14_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_4 = mask_14_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_5 = mask_14_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_6 = mask_14_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_0_7 = mask_14_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_0 = mask_14_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_1 = mask_14_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_2 = mask_14_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_3 = mask_14_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_4 = mask_14_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_5 = mask_14_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_6 = mask_14_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_1_7 = mask_14_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_0 = mask_14_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_1 = mask_14_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_2 = mask_14_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_3 = mask_14_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_4 = mask_14_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_5 = mask_14_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_6 = mask_14_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_2_7 = mask_14_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_0 = mask_14_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_1 = mask_14_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_2 = mask_14_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_3 = mask_14_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_4 = mask_14_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_5 = mask_14_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_6 = mask_14_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_3_7 = mask_14_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_0 = mask_14_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_1 = mask_14_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_2 = mask_14_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_3 = mask_14_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_4 = mask_14_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_5 = mask_14_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_6 = mask_14_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_4_7 = mask_14_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_0 = mask_14_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_1 = mask_14_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_2 = mask_14_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_3 = mask_14_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_4 = mask_14_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_5 = mask_14_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_6 = mask_14_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_5_7 = mask_14_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_0 = mask_14_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_1 = mask_14_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_2 = mask_14_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_3 = mask_14_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_4 = mask_14_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_5 = mask_14_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_6 = mask_14_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_6_7 = mask_14_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_0 = mask_14_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_1 = mask_14_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_2 = mask_14_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_3 = mask_14_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_4 = mask_14_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_5 = mask_14_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_6 = mask_14_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_14_7_7 = mask_14_7_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_0 = mask_15_0_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_1 = mask_15_0_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_2 = mask_15_0_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_3 = mask_15_0_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_4 = mask_15_0_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_5 = mask_15_0_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_6 = mask_15_0_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_0_7 = mask_15_0_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_0 = mask_15_1_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_1 = mask_15_1_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_2 = mask_15_1_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_3 = mask_15_1_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_4 = mask_15_1_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_5 = mask_15_1_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_6 = mask_15_1_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_1_7 = mask_15_1_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_0 = mask_15_2_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_1 = mask_15_2_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_2 = mask_15_2_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_3 = mask_15_2_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_4 = mask_15_2_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_5 = mask_15_2_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_6 = mask_15_2_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_2_7 = mask_15_2_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_0 = mask_15_3_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_1 = mask_15_3_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_2 = mask_15_3_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_3 = mask_15_3_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_4 = mask_15_3_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_5 = mask_15_3_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_6 = mask_15_3_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_3_7 = mask_15_3_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_0 = mask_15_4_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_1 = mask_15_4_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_2 = mask_15_4_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_3 = mask_15_4_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_4 = mask_15_4_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_5 = mask_15_4_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_6 = mask_15_4_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_4_7 = mask_15_4_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_0 = mask_15_5_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_1 = mask_15_5_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_2 = mask_15_5_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_3 = mask_15_5_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_4 = mask_15_5_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_5 = mask_15_5_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_6 = mask_15_5_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_5_7 = mask_15_5_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_0 = mask_15_6_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_1 = mask_15_6_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_2 = mask_15_6_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_3 = mask_15_6_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_4 = mask_15_6_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_5 = mask_15_6_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_6 = mask_15_6_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_6_7 = mask_15_6_7; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_0 = mask_15_7_0; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_1 = mask_15_7_1; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_2 = mask_15_7_2; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_3 = mask_15_7_3; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_4 = mask_15_7_4; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_5 = mask_15_7_5; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_6 = mask_15_7_6; // @[Sbuffer.scala 225:14]
  assign io_maskOut_15_7_7 = mask_15_7_7; // @[Sbuffer.scala 225:14]
  always @(posedge clock) begin
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_0 <= _GEN_4128;
      end
    end else begin
      data_0_0_0 <= _GEN_4128;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_1 <= _GEN_4192;
      end
    end else begin
      data_0_0_1 <= _GEN_4192;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_2 <= _GEN_4256;
      end
    end else begin
      data_0_0_2 <= _GEN_4256;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_3 <= _GEN_4320;
      end
    end else begin
      data_0_0_3 <= _GEN_4320;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_4 <= _GEN_4384;
      end
    end else begin
      data_0_0_4 <= _GEN_4384;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_5 <= _GEN_4448;
      end
    end else begin
      data_0_0_5 <= _GEN_4448;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_6 <= _GEN_4512;
      end
    end else begin
      data_0_0_6 <= _GEN_4512;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_0_7 <= _GEN_4576;
      end
    end else begin
      data_0_0_7 <= _GEN_4576;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_0 <= _GEN_4640;
      end
    end else begin
      data_0_1_0 <= _GEN_4640;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_1 <= _GEN_4704;
      end
    end else begin
      data_0_1_1 <= _GEN_4704;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_2 <= _GEN_4768;
      end
    end else begin
      data_0_1_2 <= _GEN_4768;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_3 <= _GEN_4832;
      end
    end else begin
      data_0_1_3 <= _GEN_4832;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_4 <= _GEN_4896;
      end
    end else begin
      data_0_1_4 <= _GEN_4896;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_5 <= _GEN_4960;
      end
    end else begin
      data_0_1_5 <= _GEN_4960;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_6 <= _GEN_5024;
      end
    end else begin
      data_0_1_6 <= _GEN_5024;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_1_7 <= _GEN_5088;
      end
    end else begin
      data_0_1_7 <= _GEN_5088;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_0 <= _GEN_5152;
      end
    end else begin
      data_0_2_0 <= _GEN_5152;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_1 <= _GEN_5216;
      end
    end else begin
      data_0_2_1 <= _GEN_5216;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_2 <= _GEN_5280;
      end
    end else begin
      data_0_2_2 <= _GEN_5280;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_3 <= _GEN_5344;
      end
    end else begin
      data_0_2_3 <= _GEN_5344;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_4 <= _GEN_5408;
      end
    end else begin
      data_0_2_4 <= _GEN_5408;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_5 <= _GEN_5472;
      end
    end else begin
      data_0_2_5 <= _GEN_5472;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_6 <= _GEN_5536;
      end
    end else begin
      data_0_2_6 <= _GEN_5536;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_2_7 <= _GEN_5600;
      end
    end else begin
      data_0_2_7 <= _GEN_5600;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_0 <= _GEN_5664;
      end
    end else begin
      data_0_3_0 <= _GEN_5664;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_1 <= _GEN_5728;
      end
    end else begin
      data_0_3_1 <= _GEN_5728;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_2 <= _GEN_5792;
      end
    end else begin
      data_0_3_2 <= _GEN_5792;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_3 <= _GEN_5856;
      end
    end else begin
      data_0_3_3 <= _GEN_5856;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_4 <= _GEN_5920;
      end
    end else begin
      data_0_3_4 <= _GEN_5920;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_5 <= _GEN_5984;
      end
    end else begin
      data_0_3_5 <= _GEN_5984;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_6 <= _GEN_6048;
      end
    end else begin
      data_0_3_6 <= _GEN_6048;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_3_7 <= _GEN_6112;
      end
    end else begin
      data_0_3_7 <= _GEN_6112;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_0 <= _GEN_6176;
      end
    end else begin
      data_0_4_0 <= _GEN_6176;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_1 <= _GEN_6240;
      end
    end else begin
      data_0_4_1 <= _GEN_6240;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_2 <= _GEN_6304;
      end
    end else begin
      data_0_4_2 <= _GEN_6304;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_3 <= _GEN_6368;
      end
    end else begin
      data_0_4_3 <= _GEN_6368;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_4 <= _GEN_6432;
      end
    end else begin
      data_0_4_4 <= _GEN_6432;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_5 <= _GEN_6496;
      end
    end else begin
      data_0_4_5 <= _GEN_6496;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_6 <= _GEN_6560;
      end
    end else begin
      data_0_4_6 <= _GEN_6560;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_4_7 <= _GEN_6624;
      end
    end else begin
      data_0_4_7 <= _GEN_6624;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_0 <= _GEN_6688;
      end
    end else begin
      data_0_5_0 <= _GEN_6688;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_1 <= _GEN_6752;
      end
    end else begin
      data_0_5_1 <= _GEN_6752;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_2 <= _GEN_6816;
      end
    end else begin
      data_0_5_2 <= _GEN_6816;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_3 <= _GEN_6880;
      end
    end else begin
      data_0_5_3 <= _GEN_6880;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_4 <= _GEN_6944;
      end
    end else begin
      data_0_5_4 <= _GEN_6944;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_5 <= _GEN_7008;
      end
    end else begin
      data_0_5_5 <= _GEN_7008;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_6 <= _GEN_7072;
      end
    end else begin
      data_0_5_6 <= _GEN_7072;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_5_7 <= _GEN_7136;
      end
    end else begin
      data_0_5_7 <= _GEN_7136;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_0 <= _GEN_7200;
      end
    end else begin
      data_0_6_0 <= _GEN_7200;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_1 <= _GEN_7264;
      end
    end else begin
      data_0_6_1 <= _GEN_7264;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_2 <= _GEN_7328;
      end
    end else begin
      data_0_6_2 <= _GEN_7328;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_3 <= _GEN_7392;
      end
    end else begin
      data_0_6_3 <= _GEN_7392;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_4 <= _GEN_7456;
      end
    end else begin
      data_0_6_4 <= _GEN_7456;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_5 <= _GEN_7520;
      end
    end else begin
      data_0_6_5 <= _GEN_7520;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_6 <= _GEN_7584;
      end
    end else begin
      data_0_6_6 <= _GEN_7584;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_6_7 <= _GEN_7648;
      end
    end else begin
      data_0_6_7 <= _GEN_7648;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_0 <= _GEN_7712;
      end
    end else begin
      data_0_7_0 <= _GEN_7712;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_1 <= _GEN_7776;
      end
    end else begin
      data_0_7_1 <= _GEN_7776;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_2 <= _GEN_7840;
      end
    end else begin
      data_0_7_2 <= _GEN_7840;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_3 <= _GEN_7904;
      end
    end else begin
      data_0_7_3 <= _GEN_7904;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_4 <= _GEN_7968;
      end
    end else begin
      data_0_7_4 <= _GEN_7968;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_5 <= _GEN_8032;
      end
    end else begin
      data_0_7_5 <= _GEN_8032;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_6 <= _GEN_8096;
      end
    end else begin
      data_0_7_6 <= _GEN_8096;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h0 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_0_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_0_7_7 <= _GEN_8160;
      end
    end else begin
      data_0_7_7 <= _GEN_8160;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_0 <= _GEN_4129;
      end
    end else begin
      data_1_0_0 <= _GEN_4129;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_1 <= _GEN_4193;
      end
    end else begin
      data_1_0_1 <= _GEN_4193;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_2 <= _GEN_4257;
      end
    end else begin
      data_1_0_2 <= _GEN_4257;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_3 <= _GEN_4321;
      end
    end else begin
      data_1_0_3 <= _GEN_4321;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_4 <= _GEN_4385;
      end
    end else begin
      data_1_0_4 <= _GEN_4385;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_5 <= _GEN_4449;
      end
    end else begin
      data_1_0_5 <= _GEN_4449;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_6 <= _GEN_4513;
      end
    end else begin
      data_1_0_6 <= _GEN_4513;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_0_7 <= _GEN_4577;
      end
    end else begin
      data_1_0_7 <= _GEN_4577;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_0 <= _GEN_4641;
      end
    end else begin
      data_1_1_0 <= _GEN_4641;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_1 <= _GEN_4705;
      end
    end else begin
      data_1_1_1 <= _GEN_4705;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_2 <= _GEN_4769;
      end
    end else begin
      data_1_1_2 <= _GEN_4769;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_3 <= _GEN_4833;
      end
    end else begin
      data_1_1_3 <= _GEN_4833;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_4 <= _GEN_4897;
      end
    end else begin
      data_1_1_4 <= _GEN_4897;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_5 <= _GEN_4961;
      end
    end else begin
      data_1_1_5 <= _GEN_4961;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_6 <= _GEN_5025;
      end
    end else begin
      data_1_1_6 <= _GEN_5025;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_1_7 <= _GEN_5089;
      end
    end else begin
      data_1_1_7 <= _GEN_5089;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_0 <= _GEN_5153;
      end
    end else begin
      data_1_2_0 <= _GEN_5153;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_1 <= _GEN_5217;
      end
    end else begin
      data_1_2_1 <= _GEN_5217;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_2 <= _GEN_5281;
      end
    end else begin
      data_1_2_2 <= _GEN_5281;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_3 <= _GEN_5345;
      end
    end else begin
      data_1_2_3 <= _GEN_5345;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_4 <= _GEN_5409;
      end
    end else begin
      data_1_2_4 <= _GEN_5409;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_5 <= _GEN_5473;
      end
    end else begin
      data_1_2_5 <= _GEN_5473;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_6 <= _GEN_5537;
      end
    end else begin
      data_1_2_6 <= _GEN_5537;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_2_7 <= _GEN_5601;
      end
    end else begin
      data_1_2_7 <= _GEN_5601;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_0 <= _GEN_5665;
      end
    end else begin
      data_1_3_0 <= _GEN_5665;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_1 <= _GEN_5729;
      end
    end else begin
      data_1_3_1 <= _GEN_5729;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_2 <= _GEN_5793;
      end
    end else begin
      data_1_3_2 <= _GEN_5793;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_3 <= _GEN_5857;
      end
    end else begin
      data_1_3_3 <= _GEN_5857;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_4 <= _GEN_5921;
      end
    end else begin
      data_1_3_4 <= _GEN_5921;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_5 <= _GEN_5985;
      end
    end else begin
      data_1_3_5 <= _GEN_5985;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_6 <= _GEN_6049;
      end
    end else begin
      data_1_3_6 <= _GEN_6049;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_3_7 <= _GEN_6113;
      end
    end else begin
      data_1_3_7 <= _GEN_6113;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_0 <= _GEN_6177;
      end
    end else begin
      data_1_4_0 <= _GEN_6177;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_1 <= _GEN_6241;
      end
    end else begin
      data_1_4_1 <= _GEN_6241;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_2 <= _GEN_6305;
      end
    end else begin
      data_1_4_2 <= _GEN_6305;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_3 <= _GEN_6369;
      end
    end else begin
      data_1_4_3 <= _GEN_6369;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_4 <= _GEN_6433;
      end
    end else begin
      data_1_4_4 <= _GEN_6433;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_5 <= _GEN_6497;
      end
    end else begin
      data_1_4_5 <= _GEN_6497;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_6 <= _GEN_6561;
      end
    end else begin
      data_1_4_6 <= _GEN_6561;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_4_7 <= _GEN_6625;
      end
    end else begin
      data_1_4_7 <= _GEN_6625;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_0 <= _GEN_6689;
      end
    end else begin
      data_1_5_0 <= _GEN_6689;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_1 <= _GEN_6753;
      end
    end else begin
      data_1_5_1 <= _GEN_6753;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_2 <= _GEN_6817;
      end
    end else begin
      data_1_5_2 <= _GEN_6817;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_3 <= _GEN_6881;
      end
    end else begin
      data_1_5_3 <= _GEN_6881;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_4 <= _GEN_6945;
      end
    end else begin
      data_1_5_4 <= _GEN_6945;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_5 <= _GEN_7009;
      end
    end else begin
      data_1_5_5 <= _GEN_7009;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_6 <= _GEN_7073;
      end
    end else begin
      data_1_5_6 <= _GEN_7073;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_5_7 <= _GEN_7137;
      end
    end else begin
      data_1_5_7 <= _GEN_7137;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_0 <= _GEN_7201;
      end
    end else begin
      data_1_6_0 <= _GEN_7201;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_1 <= _GEN_7265;
      end
    end else begin
      data_1_6_1 <= _GEN_7265;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_2 <= _GEN_7329;
      end
    end else begin
      data_1_6_2 <= _GEN_7329;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_3 <= _GEN_7393;
      end
    end else begin
      data_1_6_3 <= _GEN_7393;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_4 <= _GEN_7457;
      end
    end else begin
      data_1_6_4 <= _GEN_7457;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_5 <= _GEN_7521;
      end
    end else begin
      data_1_6_5 <= _GEN_7521;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_6 <= _GEN_7585;
      end
    end else begin
      data_1_6_6 <= _GEN_7585;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_6_7 <= _GEN_7649;
      end
    end else begin
      data_1_6_7 <= _GEN_7649;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_0 <= _GEN_7713;
      end
    end else begin
      data_1_7_0 <= _GEN_7713;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_1 <= _GEN_7777;
      end
    end else begin
      data_1_7_1 <= _GEN_7777;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_2 <= _GEN_7841;
      end
    end else begin
      data_1_7_2 <= _GEN_7841;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_3 <= _GEN_7905;
      end
    end else begin
      data_1_7_3 <= _GEN_7905;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_4 <= _GEN_7969;
      end
    end else begin
      data_1_7_4 <= _GEN_7969;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_5 <= _GEN_8033;
      end
    end else begin
      data_1_7_5 <= _GEN_8033;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_6 <= _GEN_8097;
      end
    end else begin
      data_1_7_6 <= _GEN_8097;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h1 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_1_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_1_7_7 <= _GEN_8161;
      end
    end else begin
      data_1_7_7 <= _GEN_8161;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_0 <= _GEN_4130;
      end
    end else begin
      data_2_0_0 <= _GEN_4130;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_1 <= _GEN_4194;
      end
    end else begin
      data_2_0_1 <= _GEN_4194;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_2 <= _GEN_4258;
      end
    end else begin
      data_2_0_2 <= _GEN_4258;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_3 <= _GEN_4322;
      end
    end else begin
      data_2_0_3 <= _GEN_4322;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_4 <= _GEN_4386;
      end
    end else begin
      data_2_0_4 <= _GEN_4386;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_5 <= _GEN_4450;
      end
    end else begin
      data_2_0_5 <= _GEN_4450;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_6 <= _GEN_4514;
      end
    end else begin
      data_2_0_6 <= _GEN_4514;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_0_7 <= _GEN_4578;
      end
    end else begin
      data_2_0_7 <= _GEN_4578;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_0 <= _GEN_4642;
      end
    end else begin
      data_2_1_0 <= _GEN_4642;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_1 <= _GEN_4706;
      end
    end else begin
      data_2_1_1 <= _GEN_4706;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_2 <= _GEN_4770;
      end
    end else begin
      data_2_1_2 <= _GEN_4770;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_3 <= _GEN_4834;
      end
    end else begin
      data_2_1_3 <= _GEN_4834;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_4 <= _GEN_4898;
      end
    end else begin
      data_2_1_4 <= _GEN_4898;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_5 <= _GEN_4962;
      end
    end else begin
      data_2_1_5 <= _GEN_4962;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_6 <= _GEN_5026;
      end
    end else begin
      data_2_1_6 <= _GEN_5026;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_1_7 <= _GEN_5090;
      end
    end else begin
      data_2_1_7 <= _GEN_5090;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_0 <= _GEN_5154;
      end
    end else begin
      data_2_2_0 <= _GEN_5154;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_1 <= _GEN_5218;
      end
    end else begin
      data_2_2_1 <= _GEN_5218;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_2 <= _GEN_5282;
      end
    end else begin
      data_2_2_2 <= _GEN_5282;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_3 <= _GEN_5346;
      end
    end else begin
      data_2_2_3 <= _GEN_5346;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_4 <= _GEN_5410;
      end
    end else begin
      data_2_2_4 <= _GEN_5410;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_5 <= _GEN_5474;
      end
    end else begin
      data_2_2_5 <= _GEN_5474;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_6 <= _GEN_5538;
      end
    end else begin
      data_2_2_6 <= _GEN_5538;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_2_7 <= _GEN_5602;
      end
    end else begin
      data_2_2_7 <= _GEN_5602;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_0 <= _GEN_5666;
      end
    end else begin
      data_2_3_0 <= _GEN_5666;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_1 <= _GEN_5730;
      end
    end else begin
      data_2_3_1 <= _GEN_5730;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_2 <= _GEN_5794;
      end
    end else begin
      data_2_3_2 <= _GEN_5794;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_3 <= _GEN_5858;
      end
    end else begin
      data_2_3_3 <= _GEN_5858;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_4 <= _GEN_5922;
      end
    end else begin
      data_2_3_4 <= _GEN_5922;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_5 <= _GEN_5986;
      end
    end else begin
      data_2_3_5 <= _GEN_5986;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_6 <= _GEN_6050;
      end
    end else begin
      data_2_3_6 <= _GEN_6050;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_3_7 <= _GEN_6114;
      end
    end else begin
      data_2_3_7 <= _GEN_6114;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_0 <= _GEN_6178;
      end
    end else begin
      data_2_4_0 <= _GEN_6178;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_1 <= _GEN_6242;
      end
    end else begin
      data_2_4_1 <= _GEN_6242;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_2 <= _GEN_6306;
      end
    end else begin
      data_2_4_2 <= _GEN_6306;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_3 <= _GEN_6370;
      end
    end else begin
      data_2_4_3 <= _GEN_6370;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_4 <= _GEN_6434;
      end
    end else begin
      data_2_4_4 <= _GEN_6434;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_5 <= _GEN_6498;
      end
    end else begin
      data_2_4_5 <= _GEN_6498;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_6 <= _GEN_6562;
      end
    end else begin
      data_2_4_6 <= _GEN_6562;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_4_7 <= _GEN_6626;
      end
    end else begin
      data_2_4_7 <= _GEN_6626;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_0 <= _GEN_6690;
      end
    end else begin
      data_2_5_0 <= _GEN_6690;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_1 <= _GEN_6754;
      end
    end else begin
      data_2_5_1 <= _GEN_6754;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_2 <= _GEN_6818;
      end
    end else begin
      data_2_5_2 <= _GEN_6818;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_3 <= _GEN_6882;
      end
    end else begin
      data_2_5_3 <= _GEN_6882;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_4 <= _GEN_6946;
      end
    end else begin
      data_2_5_4 <= _GEN_6946;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_5 <= _GEN_7010;
      end
    end else begin
      data_2_5_5 <= _GEN_7010;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_6 <= _GEN_7074;
      end
    end else begin
      data_2_5_6 <= _GEN_7074;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_5_7 <= _GEN_7138;
      end
    end else begin
      data_2_5_7 <= _GEN_7138;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_0 <= _GEN_7202;
      end
    end else begin
      data_2_6_0 <= _GEN_7202;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_1 <= _GEN_7266;
      end
    end else begin
      data_2_6_1 <= _GEN_7266;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_2 <= _GEN_7330;
      end
    end else begin
      data_2_6_2 <= _GEN_7330;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_3 <= _GEN_7394;
      end
    end else begin
      data_2_6_3 <= _GEN_7394;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_4 <= _GEN_7458;
      end
    end else begin
      data_2_6_4 <= _GEN_7458;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_5 <= _GEN_7522;
      end
    end else begin
      data_2_6_5 <= _GEN_7522;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_6 <= _GEN_7586;
      end
    end else begin
      data_2_6_6 <= _GEN_7586;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_6_7 <= _GEN_7650;
      end
    end else begin
      data_2_6_7 <= _GEN_7650;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_0 <= _GEN_7714;
      end
    end else begin
      data_2_7_0 <= _GEN_7714;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_1 <= _GEN_7778;
      end
    end else begin
      data_2_7_1 <= _GEN_7778;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_2 <= _GEN_7842;
      end
    end else begin
      data_2_7_2 <= _GEN_7842;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_3 <= _GEN_7906;
      end
    end else begin
      data_2_7_3 <= _GEN_7906;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_4 <= _GEN_7970;
      end
    end else begin
      data_2_7_4 <= _GEN_7970;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_5 <= _GEN_8034;
      end
    end else begin
      data_2_7_5 <= _GEN_8034;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_6 <= _GEN_8098;
      end
    end else begin
      data_2_7_6 <= _GEN_8098;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h2 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_2_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_2_7_7 <= _GEN_8162;
      end
    end else begin
      data_2_7_7 <= _GEN_8162;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_0 <= _GEN_4131;
      end
    end else begin
      data_3_0_0 <= _GEN_4131;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_1 <= _GEN_4195;
      end
    end else begin
      data_3_0_1 <= _GEN_4195;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_2 <= _GEN_4259;
      end
    end else begin
      data_3_0_2 <= _GEN_4259;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_3 <= _GEN_4323;
      end
    end else begin
      data_3_0_3 <= _GEN_4323;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_4 <= _GEN_4387;
      end
    end else begin
      data_3_0_4 <= _GEN_4387;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_5 <= _GEN_4451;
      end
    end else begin
      data_3_0_5 <= _GEN_4451;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_6 <= _GEN_4515;
      end
    end else begin
      data_3_0_6 <= _GEN_4515;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_0_7 <= _GEN_4579;
      end
    end else begin
      data_3_0_7 <= _GEN_4579;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_0 <= _GEN_4643;
      end
    end else begin
      data_3_1_0 <= _GEN_4643;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_1 <= _GEN_4707;
      end
    end else begin
      data_3_1_1 <= _GEN_4707;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_2 <= _GEN_4771;
      end
    end else begin
      data_3_1_2 <= _GEN_4771;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_3 <= _GEN_4835;
      end
    end else begin
      data_3_1_3 <= _GEN_4835;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_4 <= _GEN_4899;
      end
    end else begin
      data_3_1_4 <= _GEN_4899;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_5 <= _GEN_4963;
      end
    end else begin
      data_3_1_5 <= _GEN_4963;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_6 <= _GEN_5027;
      end
    end else begin
      data_3_1_6 <= _GEN_5027;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_1_7 <= _GEN_5091;
      end
    end else begin
      data_3_1_7 <= _GEN_5091;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_0 <= _GEN_5155;
      end
    end else begin
      data_3_2_0 <= _GEN_5155;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_1 <= _GEN_5219;
      end
    end else begin
      data_3_2_1 <= _GEN_5219;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_2 <= _GEN_5283;
      end
    end else begin
      data_3_2_2 <= _GEN_5283;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_3 <= _GEN_5347;
      end
    end else begin
      data_3_2_3 <= _GEN_5347;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_4 <= _GEN_5411;
      end
    end else begin
      data_3_2_4 <= _GEN_5411;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_5 <= _GEN_5475;
      end
    end else begin
      data_3_2_5 <= _GEN_5475;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_6 <= _GEN_5539;
      end
    end else begin
      data_3_2_6 <= _GEN_5539;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_2_7 <= _GEN_5603;
      end
    end else begin
      data_3_2_7 <= _GEN_5603;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_0 <= _GEN_5667;
      end
    end else begin
      data_3_3_0 <= _GEN_5667;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_1 <= _GEN_5731;
      end
    end else begin
      data_3_3_1 <= _GEN_5731;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_2 <= _GEN_5795;
      end
    end else begin
      data_3_3_2 <= _GEN_5795;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_3 <= _GEN_5859;
      end
    end else begin
      data_3_3_3 <= _GEN_5859;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_4 <= _GEN_5923;
      end
    end else begin
      data_3_3_4 <= _GEN_5923;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_5 <= _GEN_5987;
      end
    end else begin
      data_3_3_5 <= _GEN_5987;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_6 <= _GEN_6051;
      end
    end else begin
      data_3_3_6 <= _GEN_6051;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_3_7 <= _GEN_6115;
      end
    end else begin
      data_3_3_7 <= _GEN_6115;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_0 <= _GEN_6179;
      end
    end else begin
      data_3_4_0 <= _GEN_6179;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_1 <= _GEN_6243;
      end
    end else begin
      data_3_4_1 <= _GEN_6243;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_2 <= _GEN_6307;
      end
    end else begin
      data_3_4_2 <= _GEN_6307;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_3 <= _GEN_6371;
      end
    end else begin
      data_3_4_3 <= _GEN_6371;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_4 <= _GEN_6435;
      end
    end else begin
      data_3_4_4 <= _GEN_6435;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_5 <= _GEN_6499;
      end
    end else begin
      data_3_4_5 <= _GEN_6499;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_6 <= _GEN_6563;
      end
    end else begin
      data_3_4_6 <= _GEN_6563;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_4_7 <= _GEN_6627;
      end
    end else begin
      data_3_4_7 <= _GEN_6627;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_0 <= _GEN_6691;
      end
    end else begin
      data_3_5_0 <= _GEN_6691;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_1 <= _GEN_6755;
      end
    end else begin
      data_3_5_1 <= _GEN_6755;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_2 <= _GEN_6819;
      end
    end else begin
      data_3_5_2 <= _GEN_6819;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_3 <= _GEN_6883;
      end
    end else begin
      data_3_5_3 <= _GEN_6883;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_4 <= _GEN_6947;
      end
    end else begin
      data_3_5_4 <= _GEN_6947;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_5 <= _GEN_7011;
      end
    end else begin
      data_3_5_5 <= _GEN_7011;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_6 <= _GEN_7075;
      end
    end else begin
      data_3_5_6 <= _GEN_7075;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_5_7 <= _GEN_7139;
      end
    end else begin
      data_3_5_7 <= _GEN_7139;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_0 <= _GEN_7203;
      end
    end else begin
      data_3_6_0 <= _GEN_7203;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_1 <= _GEN_7267;
      end
    end else begin
      data_3_6_1 <= _GEN_7267;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_2 <= _GEN_7331;
      end
    end else begin
      data_3_6_2 <= _GEN_7331;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_3 <= _GEN_7395;
      end
    end else begin
      data_3_6_3 <= _GEN_7395;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_4 <= _GEN_7459;
      end
    end else begin
      data_3_6_4 <= _GEN_7459;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_5 <= _GEN_7523;
      end
    end else begin
      data_3_6_5 <= _GEN_7523;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_6 <= _GEN_7587;
      end
    end else begin
      data_3_6_6 <= _GEN_7587;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_6_7 <= _GEN_7651;
      end
    end else begin
      data_3_6_7 <= _GEN_7651;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_0 <= _GEN_7715;
      end
    end else begin
      data_3_7_0 <= _GEN_7715;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_1 <= _GEN_7779;
      end
    end else begin
      data_3_7_1 <= _GEN_7779;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_2 <= _GEN_7843;
      end
    end else begin
      data_3_7_2 <= _GEN_7843;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_3 <= _GEN_7907;
      end
    end else begin
      data_3_7_3 <= _GEN_7907;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_4 <= _GEN_7971;
      end
    end else begin
      data_3_7_4 <= _GEN_7971;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_5 <= _GEN_8035;
      end
    end else begin
      data_3_7_5 <= _GEN_8035;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_6 <= _GEN_8099;
      end
    end else begin
      data_3_7_6 <= _GEN_8099;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h3 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_3_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_3_7_7 <= _GEN_8163;
      end
    end else begin
      data_3_7_7 <= _GEN_8163;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_0 <= _GEN_4132;
      end
    end else begin
      data_4_0_0 <= _GEN_4132;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_1 <= _GEN_4196;
      end
    end else begin
      data_4_0_1 <= _GEN_4196;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_2 <= _GEN_4260;
      end
    end else begin
      data_4_0_2 <= _GEN_4260;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_3 <= _GEN_4324;
      end
    end else begin
      data_4_0_3 <= _GEN_4324;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_4 <= _GEN_4388;
      end
    end else begin
      data_4_0_4 <= _GEN_4388;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_5 <= _GEN_4452;
      end
    end else begin
      data_4_0_5 <= _GEN_4452;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_6 <= _GEN_4516;
      end
    end else begin
      data_4_0_6 <= _GEN_4516;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_0_7 <= _GEN_4580;
      end
    end else begin
      data_4_0_7 <= _GEN_4580;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_0 <= _GEN_4644;
      end
    end else begin
      data_4_1_0 <= _GEN_4644;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_1 <= _GEN_4708;
      end
    end else begin
      data_4_1_1 <= _GEN_4708;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_2 <= _GEN_4772;
      end
    end else begin
      data_4_1_2 <= _GEN_4772;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_3 <= _GEN_4836;
      end
    end else begin
      data_4_1_3 <= _GEN_4836;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_4 <= _GEN_4900;
      end
    end else begin
      data_4_1_4 <= _GEN_4900;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_5 <= _GEN_4964;
      end
    end else begin
      data_4_1_5 <= _GEN_4964;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_6 <= _GEN_5028;
      end
    end else begin
      data_4_1_6 <= _GEN_5028;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_1_7 <= _GEN_5092;
      end
    end else begin
      data_4_1_7 <= _GEN_5092;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_0 <= _GEN_5156;
      end
    end else begin
      data_4_2_0 <= _GEN_5156;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_1 <= _GEN_5220;
      end
    end else begin
      data_4_2_1 <= _GEN_5220;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_2 <= _GEN_5284;
      end
    end else begin
      data_4_2_2 <= _GEN_5284;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_3 <= _GEN_5348;
      end
    end else begin
      data_4_2_3 <= _GEN_5348;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_4 <= _GEN_5412;
      end
    end else begin
      data_4_2_4 <= _GEN_5412;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_5 <= _GEN_5476;
      end
    end else begin
      data_4_2_5 <= _GEN_5476;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_6 <= _GEN_5540;
      end
    end else begin
      data_4_2_6 <= _GEN_5540;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_2_7 <= _GEN_5604;
      end
    end else begin
      data_4_2_7 <= _GEN_5604;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_0 <= _GEN_5668;
      end
    end else begin
      data_4_3_0 <= _GEN_5668;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_1 <= _GEN_5732;
      end
    end else begin
      data_4_3_1 <= _GEN_5732;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_2 <= _GEN_5796;
      end
    end else begin
      data_4_3_2 <= _GEN_5796;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_3 <= _GEN_5860;
      end
    end else begin
      data_4_3_3 <= _GEN_5860;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_4 <= _GEN_5924;
      end
    end else begin
      data_4_3_4 <= _GEN_5924;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_5 <= _GEN_5988;
      end
    end else begin
      data_4_3_5 <= _GEN_5988;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_6 <= _GEN_6052;
      end
    end else begin
      data_4_3_6 <= _GEN_6052;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_3_7 <= _GEN_6116;
      end
    end else begin
      data_4_3_7 <= _GEN_6116;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_0 <= _GEN_6180;
      end
    end else begin
      data_4_4_0 <= _GEN_6180;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_1 <= _GEN_6244;
      end
    end else begin
      data_4_4_1 <= _GEN_6244;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_2 <= _GEN_6308;
      end
    end else begin
      data_4_4_2 <= _GEN_6308;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_3 <= _GEN_6372;
      end
    end else begin
      data_4_4_3 <= _GEN_6372;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_4 <= _GEN_6436;
      end
    end else begin
      data_4_4_4 <= _GEN_6436;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_5 <= _GEN_6500;
      end
    end else begin
      data_4_4_5 <= _GEN_6500;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_6 <= _GEN_6564;
      end
    end else begin
      data_4_4_6 <= _GEN_6564;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_4_7 <= _GEN_6628;
      end
    end else begin
      data_4_4_7 <= _GEN_6628;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_0 <= _GEN_6692;
      end
    end else begin
      data_4_5_0 <= _GEN_6692;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_1 <= _GEN_6756;
      end
    end else begin
      data_4_5_1 <= _GEN_6756;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_2 <= _GEN_6820;
      end
    end else begin
      data_4_5_2 <= _GEN_6820;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_3 <= _GEN_6884;
      end
    end else begin
      data_4_5_3 <= _GEN_6884;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_4 <= _GEN_6948;
      end
    end else begin
      data_4_5_4 <= _GEN_6948;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_5 <= _GEN_7012;
      end
    end else begin
      data_4_5_5 <= _GEN_7012;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_6 <= _GEN_7076;
      end
    end else begin
      data_4_5_6 <= _GEN_7076;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_5_7 <= _GEN_7140;
      end
    end else begin
      data_4_5_7 <= _GEN_7140;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_0 <= _GEN_7204;
      end
    end else begin
      data_4_6_0 <= _GEN_7204;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_1 <= _GEN_7268;
      end
    end else begin
      data_4_6_1 <= _GEN_7268;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_2 <= _GEN_7332;
      end
    end else begin
      data_4_6_2 <= _GEN_7332;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_3 <= _GEN_7396;
      end
    end else begin
      data_4_6_3 <= _GEN_7396;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_4 <= _GEN_7460;
      end
    end else begin
      data_4_6_4 <= _GEN_7460;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_5 <= _GEN_7524;
      end
    end else begin
      data_4_6_5 <= _GEN_7524;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_6 <= _GEN_7588;
      end
    end else begin
      data_4_6_6 <= _GEN_7588;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_6_7 <= _GEN_7652;
      end
    end else begin
      data_4_6_7 <= _GEN_7652;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_0 <= _GEN_7716;
      end
    end else begin
      data_4_7_0 <= _GEN_7716;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_1 <= _GEN_7780;
      end
    end else begin
      data_4_7_1 <= _GEN_7780;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_2 <= _GEN_7844;
      end
    end else begin
      data_4_7_2 <= _GEN_7844;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_3 <= _GEN_7908;
      end
    end else begin
      data_4_7_3 <= _GEN_7908;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_4 <= _GEN_7972;
      end
    end else begin
      data_4_7_4 <= _GEN_7972;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_5 <= _GEN_8036;
      end
    end else begin
      data_4_7_5 <= _GEN_8036;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_6 <= _GEN_8100;
      end
    end else begin
      data_4_7_6 <= _GEN_8100;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h4 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_4_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_4_7_7 <= _GEN_8164;
      end
    end else begin
      data_4_7_7 <= _GEN_8164;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_0 <= _GEN_4133;
      end
    end else begin
      data_5_0_0 <= _GEN_4133;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_1 <= _GEN_4197;
      end
    end else begin
      data_5_0_1 <= _GEN_4197;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_2 <= _GEN_4261;
      end
    end else begin
      data_5_0_2 <= _GEN_4261;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_3 <= _GEN_4325;
      end
    end else begin
      data_5_0_3 <= _GEN_4325;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_4 <= _GEN_4389;
      end
    end else begin
      data_5_0_4 <= _GEN_4389;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_5 <= _GEN_4453;
      end
    end else begin
      data_5_0_5 <= _GEN_4453;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_6 <= _GEN_4517;
      end
    end else begin
      data_5_0_6 <= _GEN_4517;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_0_7 <= _GEN_4581;
      end
    end else begin
      data_5_0_7 <= _GEN_4581;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_0 <= _GEN_4645;
      end
    end else begin
      data_5_1_0 <= _GEN_4645;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_1 <= _GEN_4709;
      end
    end else begin
      data_5_1_1 <= _GEN_4709;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_2 <= _GEN_4773;
      end
    end else begin
      data_5_1_2 <= _GEN_4773;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_3 <= _GEN_4837;
      end
    end else begin
      data_5_1_3 <= _GEN_4837;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_4 <= _GEN_4901;
      end
    end else begin
      data_5_1_4 <= _GEN_4901;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_5 <= _GEN_4965;
      end
    end else begin
      data_5_1_5 <= _GEN_4965;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_6 <= _GEN_5029;
      end
    end else begin
      data_5_1_6 <= _GEN_5029;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_1_7 <= _GEN_5093;
      end
    end else begin
      data_5_1_7 <= _GEN_5093;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_0 <= _GEN_5157;
      end
    end else begin
      data_5_2_0 <= _GEN_5157;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_1 <= _GEN_5221;
      end
    end else begin
      data_5_2_1 <= _GEN_5221;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_2 <= _GEN_5285;
      end
    end else begin
      data_5_2_2 <= _GEN_5285;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_3 <= _GEN_5349;
      end
    end else begin
      data_5_2_3 <= _GEN_5349;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_4 <= _GEN_5413;
      end
    end else begin
      data_5_2_4 <= _GEN_5413;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_5 <= _GEN_5477;
      end
    end else begin
      data_5_2_5 <= _GEN_5477;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_6 <= _GEN_5541;
      end
    end else begin
      data_5_2_6 <= _GEN_5541;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_2_7 <= _GEN_5605;
      end
    end else begin
      data_5_2_7 <= _GEN_5605;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_0 <= _GEN_5669;
      end
    end else begin
      data_5_3_0 <= _GEN_5669;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_1 <= _GEN_5733;
      end
    end else begin
      data_5_3_1 <= _GEN_5733;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_2 <= _GEN_5797;
      end
    end else begin
      data_5_3_2 <= _GEN_5797;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_3 <= _GEN_5861;
      end
    end else begin
      data_5_3_3 <= _GEN_5861;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_4 <= _GEN_5925;
      end
    end else begin
      data_5_3_4 <= _GEN_5925;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_5 <= _GEN_5989;
      end
    end else begin
      data_5_3_5 <= _GEN_5989;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_6 <= _GEN_6053;
      end
    end else begin
      data_5_3_6 <= _GEN_6053;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_3_7 <= _GEN_6117;
      end
    end else begin
      data_5_3_7 <= _GEN_6117;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_0 <= _GEN_6181;
      end
    end else begin
      data_5_4_0 <= _GEN_6181;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_1 <= _GEN_6245;
      end
    end else begin
      data_5_4_1 <= _GEN_6245;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_2 <= _GEN_6309;
      end
    end else begin
      data_5_4_2 <= _GEN_6309;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_3 <= _GEN_6373;
      end
    end else begin
      data_5_4_3 <= _GEN_6373;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_4 <= _GEN_6437;
      end
    end else begin
      data_5_4_4 <= _GEN_6437;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_5 <= _GEN_6501;
      end
    end else begin
      data_5_4_5 <= _GEN_6501;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_6 <= _GEN_6565;
      end
    end else begin
      data_5_4_6 <= _GEN_6565;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_4_7 <= _GEN_6629;
      end
    end else begin
      data_5_4_7 <= _GEN_6629;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_0 <= _GEN_6693;
      end
    end else begin
      data_5_5_0 <= _GEN_6693;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_1 <= _GEN_6757;
      end
    end else begin
      data_5_5_1 <= _GEN_6757;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_2 <= _GEN_6821;
      end
    end else begin
      data_5_5_2 <= _GEN_6821;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_3 <= _GEN_6885;
      end
    end else begin
      data_5_5_3 <= _GEN_6885;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_4 <= _GEN_6949;
      end
    end else begin
      data_5_5_4 <= _GEN_6949;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_5 <= _GEN_7013;
      end
    end else begin
      data_5_5_5 <= _GEN_7013;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_6 <= _GEN_7077;
      end
    end else begin
      data_5_5_6 <= _GEN_7077;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_5_7 <= _GEN_7141;
      end
    end else begin
      data_5_5_7 <= _GEN_7141;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_0 <= _GEN_7205;
      end
    end else begin
      data_5_6_0 <= _GEN_7205;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_1 <= _GEN_7269;
      end
    end else begin
      data_5_6_1 <= _GEN_7269;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_2 <= _GEN_7333;
      end
    end else begin
      data_5_6_2 <= _GEN_7333;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_3 <= _GEN_7397;
      end
    end else begin
      data_5_6_3 <= _GEN_7397;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_4 <= _GEN_7461;
      end
    end else begin
      data_5_6_4 <= _GEN_7461;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_5 <= _GEN_7525;
      end
    end else begin
      data_5_6_5 <= _GEN_7525;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_6 <= _GEN_7589;
      end
    end else begin
      data_5_6_6 <= _GEN_7589;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_6_7 <= _GEN_7653;
      end
    end else begin
      data_5_6_7 <= _GEN_7653;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_0 <= _GEN_7717;
      end
    end else begin
      data_5_7_0 <= _GEN_7717;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_1 <= _GEN_7781;
      end
    end else begin
      data_5_7_1 <= _GEN_7781;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_2 <= _GEN_7845;
      end
    end else begin
      data_5_7_2 <= _GEN_7845;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_3 <= _GEN_7909;
      end
    end else begin
      data_5_7_3 <= _GEN_7909;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_4 <= _GEN_7973;
      end
    end else begin
      data_5_7_4 <= _GEN_7973;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_5 <= _GEN_8037;
      end
    end else begin
      data_5_7_5 <= _GEN_8037;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_6 <= _GEN_8101;
      end
    end else begin
      data_5_7_6 <= _GEN_8101;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h5 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_5_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_5_7_7 <= _GEN_8165;
      end
    end else begin
      data_5_7_7 <= _GEN_8165;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_0 <= _GEN_4134;
      end
    end else begin
      data_6_0_0 <= _GEN_4134;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_1 <= _GEN_4198;
      end
    end else begin
      data_6_0_1 <= _GEN_4198;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_2 <= _GEN_4262;
      end
    end else begin
      data_6_0_2 <= _GEN_4262;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_3 <= _GEN_4326;
      end
    end else begin
      data_6_0_3 <= _GEN_4326;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_4 <= _GEN_4390;
      end
    end else begin
      data_6_0_4 <= _GEN_4390;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_5 <= _GEN_4454;
      end
    end else begin
      data_6_0_5 <= _GEN_4454;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_6 <= _GEN_4518;
      end
    end else begin
      data_6_0_6 <= _GEN_4518;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_0_7 <= _GEN_4582;
      end
    end else begin
      data_6_0_7 <= _GEN_4582;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_0 <= _GEN_4646;
      end
    end else begin
      data_6_1_0 <= _GEN_4646;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_1 <= _GEN_4710;
      end
    end else begin
      data_6_1_1 <= _GEN_4710;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_2 <= _GEN_4774;
      end
    end else begin
      data_6_1_2 <= _GEN_4774;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_3 <= _GEN_4838;
      end
    end else begin
      data_6_1_3 <= _GEN_4838;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_4 <= _GEN_4902;
      end
    end else begin
      data_6_1_4 <= _GEN_4902;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_5 <= _GEN_4966;
      end
    end else begin
      data_6_1_5 <= _GEN_4966;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_6 <= _GEN_5030;
      end
    end else begin
      data_6_1_6 <= _GEN_5030;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_1_7 <= _GEN_5094;
      end
    end else begin
      data_6_1_7 <= _GEN_5094;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_0 <= _GEN_5158;
      end
    end else begin
      data_6_2_0 <= _GEN_5158;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_1 <= _GEN_5222;
      end
    end else begin
      data_6_2_1 <= _GEN_5222;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_2 <= _GEN_5286;
      end
    end else begin
      data_6_2_2 <= _GEN_5286;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_3 <= _GEN_5350;
      end
    end else begin
      data_6_2_3 <= _GEN_5350;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_4 <= _GEN_5414;
      end
    end else begin
      data_6_2_4 <= _GEN_5414;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_5 <= _GEN_5478;
      end
    end else begin
      data_6_2_5 <= _GEN_5478;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_6 <= _GEN_5542;
      end
    end else begin
      data_6_2_6 <= _GEN_5542;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_2_7 <= _GEN_5606;
      end
    end else begin
      data_6_2_7 <= _GEN_5606;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_0 <= _GEN_5670;
      end
    end else begin
      data_6_3_0 <= _GEN_5670;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_1 <= _GEN_5734;
      end
    end else begin
      data_6_3_1 <= _GEN_5734;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_2 <= _GEN_5798;
      end
    end else begin
      data_6_3_2 <= _GEN_5798;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_3 <= _GEN_5862;
      end
    end else begin
      data_6_3_3 <= _GEN_5862;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_4 <= _GEN_5926;
      end
    end else begin
      data_6_3_4 <= _GEN_5926;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_5 <= _GEN_5990;
      end
    end else begin
      data_6_3_5 <= _GEN_5990;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_6 <= _GEN_6054;
      end
    end else begin
      data_6_3_6 <= _GEN_6054;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_3_7 <= _GEN_6118;
      end
    end else begin
      data_6_3_7 <= _GEN_6118;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_0 <= _GEN_6182;
      end
    end else begin
      data_6_4_0 <= _GEN_6182;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_1 <= _GEN_6246;
      end
    end else begin
      data_6_4_1 <= _GEN_6246;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_2 <= _GEN_6310;
      end
    end else begin
      data_6_4_2 <= _GEN_6310;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_3 <= _GEN_6374;
      end
    end else begin
      data_6_4_3 <= _GEN_6374;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_4 <= _GEN_6438;
      end
    end else begin
      data_6_4_4 <= _GEN_6438;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_5 <= _GEN_6502;
      end
    end else begin
      data_6_4_5 <= _GEN_6502;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_6 <= _GEN_6566;
      end
    end else begin
      data_6_4_6 <= _GEN_6566;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_4_7 <= _GEN_6630;
      end
    end else begin
      data_6_4_7 <= _GEN_6630;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_0 <= _GEN_6694;
      end
    end else begin
      data_6_5_0 <= _GEN_6694;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_1 <= _GEN_6758;
      end
    end else begin
      data_6_5_1 <= _GEN_6758;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_2 <= _GEN_6822;
      end
    end else begin
      data_6_5_2 <= _GEN_6822;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_3 <= _GEN_6886;
      end
    end else begin
      data_6_5_3 <= _GEN_6886;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_4 <= _GEN_6950;
      end
    end else begin
      data_6_5_4 <= _GEN_6950;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_5 <= _GEN_7014;
      end
    end else begin
      data_6_5_5 <= _GEN_7014;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_6 <= _GEN_7078;
      end
    end else begin
      data_6_5_6 <= _GEN_7078;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_5_7 <= _GEN_7142;
      end
    end else begin
      data_6_5_7 <= _GEN_7142;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_0 <= _GEN_7206;
      end
    end else begin
      data_6_6_0 <= _GEN_7206;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_1 <= _GEN_7270;
      end
    end else begin
      data_6_6_1 <= _GEN_7270;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_2 <= _GEN_7334;
      end
    end else begin
      data_6_6_2 <= _GEN_7334;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_3 <= _GEN_7398;
      end
    end else begin
      data_6_6_3 <= _GEN_7398;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_4 <= _GEN_7462;
      end
    end else begin
      data_6_6_4 <= _GEN_7462;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_5 <= _GEN_7526;
      end
    end else begin
      data_6_6_5 <= _GEN_7526;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_6 <= _GEN_7590;
      end
    end else begin
      data_6_6_6 <= _GEN_7590;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_6_7 <= _GEN_7654;
      end
    end else begin
      data_6_6_7 <= _GEN_7654;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_0 <= _GEN_7718;
      end
    end else begin
      data_6_7_0 <= _GEN_7718;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_1 <= _GEN_7782;
      end
    end else begin
      data_6_7_1 <= _GEN_7782;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_2 <= _GEN_7846;
      end
    end else begin
      data_6_7_2 <= _GEN_7846;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_3 <= _GEN_7910;
      end
    end else begin
      data_6_7_3 <= _GEN_7910;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_4 <= _GEN_7974;
      end
    end else begin
      data_6_7_4 <= _GEN_7974;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_5 <= _GEN_8038;
      end
    end else begin
      data_6_7_5 <= _GEN_8038;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_6 <= _GEN_8102;
      end
    end else begin
      data_6_7_6 <= _GEN_8102;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h6 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_6_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_6_7_7 <= _GEN_8166;
      end
    end else begin
      data_6_7_7 <= _GEN_8166;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_0 <= _GEN_4135;
      end
    end else begin
      data_7_0_0 <= _GEN_4135;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_1 <= _GEN_4199;
      end
    end else begin
      data_7_0_1 <= _GEN_4199;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_2 <= _GEN_4263;
      end
    end else begin
      data_7_0_2 <= _GEN_4263;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_3 <= _GEN_4327;
      end
    end else begin
      data_7_0_3 <= _GEN_4327;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_4 <= _GEN_4391;
      end
    end else begin
      data_7_0_4 <= _GEN_4391;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_5 <= _GEN_4455;
      end
    end else begin
      data_7_0_5 <= _GEN_4455;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_6 <= _GEN_4519;
      end
    end else begin
      data_7_0_6 <= _GEN_4519;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_0_7 <= _GEN_4583;
      end
    end else begin
      data_7_0_7 <= _GEN_4583;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_0 <= _GEN_4647;
      end
    end else begin
      data_7_1_0 <= _GEN_4647;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_1 <= _GEN_4711;
      end
    end else begin
      data_7_1_1 <= _GEN_4711;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_2 <= _GEN_4775;
      end
    end else begin
      data_7_1_2 <= _GEN_4775;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_3 <= _GEN_4839;
      end
    end else begin
      data_7_1_3 <= _GEN_4839;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_4 <= _GEN_4903;
      end
    end else begin
      data_7_1_4 <= _GEN_4903;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_5 <= _GEN_4967;
      end
    end else begin
      data_7_1_5 <= _GEN_4967;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_6 <= _GEN_5031;
      end
    end else begin
      data_7_1_6 <= _GEN_5031;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_1_7 <= _GEN_5095;
      end
    end else begin
      data_7_1_7 <= _GEN_5095;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_0 <= _GEN_5159;
      end
    end else begin
      data_7_2_0 <= _GEN_5159;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_1 <= _GEN_5223;
      end
    end else begin
      data_7_2_1 <= _GEN_5223;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_2 <= _GEN_5287;
      end
    end else begin
      data_7_2_2 <= _GEN_5287;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_3 <= _GEN_5351;
      end
    end else begin
      data_7_2_3 <= _GEN_5351;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_4 <= _GEN_5415;
      end
    end else begin
      data_7_2_4 <= _GEN_5415;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_5 <= _GEN_5479;
      end
    end else begin
      data_7_2_5 <= _GEN_5479;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_6 <= _GEN_5543;
      end
    end else begin
      data_7_2_6 <= _GEN_5543;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_2_7 <= _GEN_5607;
      end
    end else begin
      data_7_2_7 <= _GEN_5607;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_0 <= _GEN_5671;
      end
    end else begin
      data_7_3_0 <= _GEN_5671;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_1 <= _GEN_5735;
      end
    end else begin
      data_7_3_1 <= _GEN_5735;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_2 <= _GEN_5799;
      end
    end else begin
      data_7_3_2 <= _GEN_5799;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_3 <= _GEN_5863;
      end
    end else begin
      data_7_3_3 <= _GEN_5863;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_4 <= _GEN_5927;
      end
    end else begin
      data_7_3_4 <= _GEN_5927;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_5 <= _GEN_5991;
      end
    end else begin
      data_7_3_5 <= _GEN_5991;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_6 <= _GEN_6055;
      end
    end else begin
      data_7_3_6 <= _GEN_6055;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_3_7 <= _GEN_6119;
      end
    end else begin
      data_7_3_7 <= _GEN_6119;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_0 <= _GEN_6183;
      end
    end else begin
      data_7_4_0 <= _GEN_6183;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_1 <= _GEN_6247;
      end
    end else begin
      data_7_4_1 <= _GEN_6247;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_2 <= _GEN_6311;
      end
    end else begin
      data_7_4_2 <= _GEN_6311;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_3 <= _GEN_6375;
      end
    end else begin
      data_7_4_3 <= _GEN_6375;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_4 <= _GEN_6439;
      end
    end else begin
      data_7_4_4 <= _GEN_6439;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_5 <= _GEN_6503;
      end
    end else begin
      data_7_4_5 <= _GEN_6503;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_6 <= _GEN_6567;
      end
    end else begin
      data_7_4_6 <= _GEN_6567;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_4_7 <= _GEN_6631;
      end
    end else begin
      data_7_4_7 <= _GEN_6631;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_0 <= _GEN_6695;
      end
    end else begin
      data_7_5_0 <= _GEN_6695;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_1 <= _GEN_6759;
      end
    end else begin
      data_7_5_1 <= _GEN_6759;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_2 <= _GEN_6823;
      end
    end else begin
      data_7_5_2 <= _GEN_6823;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_3 <= _GEN_6887;
      end
    end else begin
      data_7_5_3 <= _GEN_6887;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_4 <= _GEN_6951;
      end
    end else begin
      data_7_5_4 <= _GEN_6951;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_5 <= _GEN_7015;
      end
    end else begin
      data_7_5_5 <= _GEN_7015;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_6 <= _GEN_7079;
      end
    end else begin
      data_7_5_6 <= _GEN_7079;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_5_7 <= _GEN_7143;
      end
    end else begin
      data_7_5_7 <= _GEN_7143;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_0 <= _GEN_7207;
      end
    end else begin
      data_7_6_0 <= _GEN_7207;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_1 <= _GEN_7271;
      end
    end else begin
      data_7_6_1 <= _GEN_7271;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_2 <= _GEN_7335;
      end
    end else begin
      data_7_6_2 <= _GEN_7335;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_3 <= _GEN_7399;
      end
    end else begin
      data_7_6_3 <= _GEN_7399;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_4 <= _GEN_7463;
      end
    end else begin
      data_7_6_4 <= _GEN_7463;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_5 <= _GEN_7527;
      end
    end else begin
      data_7_6_5 <= _GEN_7527;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_6 <= _GEN_7591;
      end
    end else begin
      data_7_6_6 <= _GEN_7591;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_6_7 <= _GEN_7655;
      end
    end else begin
      data_7_6_7 <= _GEN_7655;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_0 <= _GEN_7719;
      end
    end else begin
      data_7_7_0 <= _GEN_7719;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_1 <= _GEN_7783;
      end
    end else begin
      data_7_7_1 <= _GEN_7783;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_2 <= _GEN_7847;
      end
    end else begin
      data_7_7_2 <= _GEN_7847;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_3 <= _GEN_7911;
      end
    end else begin
      data_7_7_3 <= _GEN_7911;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_4 <= _GEN_7975;
      end
    end else begin
      data_7_7_4 <= _GEN_7975;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_5 <= _GEN_8039;
      end
    end else begin
      data_7_7_5 <= _GEN_8039;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_6 <= _GEN_8103;
      end
    end else begin
      data_7_7_6 <= _GEN_8103;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h7 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_7_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_7_7_7 <= _GEN_8167;
      end
    end else begin
      data_7_7_7 <= _GEN_8167;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_0 <= _GEN_4136;
      end
    end else begin
      data_8_0_0 <= _GEN_4136;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_1 <= _GEN_4200;
      end
    end else begin
      data_8_0_1 <= _GEN_4200;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_2 <= _GEN_4264;
      end
    end else begin
      data_8_0_2 <= _GEN_4264;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_3 <= _GEN_4328;
      end
    end else begin
      data_8_0_3 <= _GEN_4328;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_4 <= _GEN_4392;
      end
    end else begin
      data_8_0_4 <= _GEN_4392;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_5 <= _GEN_4456;
      end
    end else begin
      data_8_0_5 <= _GEN_4456;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_6 <= _GEN_4520;
      end
    end else begin
      data_8_0_6 <= _GEN_4520;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_0_7 <= _GEN_4584;
      end
    end else begin
      data_8_0_7 <= _GEN_4584;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_0 <= _GEN_4648;
      end
    end else begin
      data_8_1_0 <= _GEN_4648;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_1 <= _GEN_4712;
      end
    end else begin
      data_8_1_1 <= _GEN_4712;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_2 <= _GEN_4776;
      end
    end else begin
      data_8_1_2 <= _GEN_4776;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_3 <= _GEN_4840;
      end
    end else begin
      data_8_1_3 <= _GEN_4840;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_4 <= _GEN_4904;
      end
    end else begin
      data_8_1_4 <= _GEN_4904;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_5 <= _GEN_4968;
      end
    end else begin
      data_8_1_5 <= _GEN_4968;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_6 <= _GEN_5032;
      end
    end else begin
      data_8_1_6 <= _GEN_5032;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_1_7 <= _GEN_5096;
      end
    end else begin
      data_8_1_7 <= _GEN_5096;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_0 <= _GEN_5160;
      end
    end else begin
      data_8_2_0 <= _GEN_5160;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_1 <= _GEN_5224;
      end
    end else begin
      data_8_2_1 <= _GEN_5224;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_2 <= _GEN_5288;
      end
    end else begin
      data_8_2_2 <= _GEN_5288;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_3 <= _GEN_5352;
      end
    end else begin
      data_8_2_3 <= _GEN_5352;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_4 <= _GEN_5416;
      end
    end else begin
      data_8_2_4 <= _GEN_5416;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_5 <= _GEN_5480;
      end
    end else begin
      data_8_2_5 <= _GEN_5480;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_6 <= _GEN_5544;
      end
    end else begin
      data_8_2_6 <= _GEN_5544;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_2_7 <= _GEN_5608;
      end
    end else begin
      data_8_2_7 <= _GEN_5608;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_0 <= _GEN_5672;
      end
    end else begin
      data_8_3_0 <= _GEN_5672;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_1 <= _GEN_5736;
      end
    end else begin
      data_8_3_1 <= _GEN_5736;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_2 <= _GEN_5800;
      end
    end else begin
      data_8_3_2 <= _GEN_5800;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_3 <= _GEN_5864;
      end
    end else begin
      data_8_3_3 <= _GEN_5864;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_4 <= _GEN_5928;
      end
    end else begin
      data_8_3_4 <= _GEN_5928;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_5 <= _GEN_5992;
      end
    end else begin
      data_8_3_5 <= _GEN_5992;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_6 <= _GEN_6056;
      end
    end else begin
      data_8_3_6 <= _GEN_6056;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_3_7 <= _GEN_6120;
      end
    end else begin
      data_8_3_7 <= _GEN_6120;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_0 <= _GEN_6184;
      end
    end else begin
      data_8_4_0 <= _GEN_6184;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_1 <= _GEN_6248;
      end
    end else begin
      data_8_4_1 <= _GEN_6248;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_2 <= _GEN_6312;
      end
    end else begin
      data_8_4_2 <= _GEN_6312;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_3 <= _GEN_6376;
      end
    end else begin
      data_8_4_3 <= _GEN_6376;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_4 <= _GEN_6440;
      end
    end else begin
      data_8_4_4 <= _GEN_6440;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_5 <= _GEN_6504;
      end
    end else begin
      data_8_4_5 <= _GEN_6504;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_6 <= _GEN_6568;
      end
    end else begin
      data_8_4_6 <= _GEN_6568;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_4_7 <= _GEN_6632;
      end
    end else begin
      data_8_4_7 <= _GEN_6632;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_0 <= _GEN_6696;
      end
    end else begin
      data_8_5_0 <= _GEN_6696;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_1 <= _GEN_6760;
      end
    end else begin
      data_8_5_1 <= _GEN_6760;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_2 <= _GEN_6824;
      end
    end else begin
      data_8_5_2 <= _GEN_6824;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_3 <= _GEN_6888;
      end
    end else begin
      data_8_5_3 <= _GEN_6888;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_4 <= _GEN_6952;
      end
    end else begin
      data_8_5_4 <= _GEN_6952;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_5 <= _GEN_7016;
      end
    end else begin
      data_8_5_5 <= _GEN_7016;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_6 <= _GEN_7080;
      end
    end else begin
      data_8_5_6 <= _GEN_7080;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_5_7 <= _GEN_7144;
      end
    end else begin
      data_8_5_7 <= _GEN_7144;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_0 <= _GEN_7208;
      end
    end else begin
      data_8_6_0 <= _GEN_7208;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_1 <= _GEN_7272;
      end
    end else begin
      data_8_6_1 <= _GEN_7272;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_2 <= _GEN_7336;
      end
    end else begin
      data_8_6_2 <= _GEN_7336;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_3 <= _GEN_7400;
      end
    end else begin
      data_8_6_3 <= _GEN_7400;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_4 <= _GEN_7464;
      end
    end else begin
      data_8_6_4 <= _GEN_7464;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_5 <= _GEN_7528;
      end
    end else begin
      data_8_6_5 <= _GEN_7528;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_6 <= _GEN_7592;
      end
    end else begin
      data_8_6_6 <= _GEN_7592;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_6_7 <= _GEN_7656;
      end
    end else begin
      data_8_6_7 <= _GEN_7656;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_0 <= _GEN_7720;
      end
    end else begin
      data_8_7_0 <= _GEN_7720;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_1 <= _GEN_7784;
      end
    end else begin
      data_8_7_1 <= _GEN_7784;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_2 <= _GEN_7848;
      end
    end else begin
      data_8_7_2 <= _GEN_7848;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_3 <= _GEN_7912;
      end
    end else begin
      data_8_7_3 <= _GEN_7912;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_4 <= _GEN_7976;
      end
    end else begin
      data_8_7_4 <= _GEN_7976;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_5 <= _GEN_8040;
      end
    end else begin
      data_8_7_5 <= _GEN_8040;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_6 <= _GEN_8104;
      end
    end else begin
      data_8_7_6 <= _GEN_8104;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h8 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_8_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_8_7_7 <= _GEN_8168;
      end
    end else begin
      data_8_7_7 <= _GEN_8168;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_0 <= _GEN_4137;
      end
    end else begin
      data_9_0_0 <= _GEN_4137;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_1 <= _GEN_4201;
      end
    end else begin
      data_9_0_1 <= _GEN_4201;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_2 <= _GEN_4265;
      end
    end else begin
      data_9_0_2 <= _GEN_4265;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_3 <= _GEN_4329;
      end
    end else begin
      data_9_0_3 <= _GEN_4329;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_4 <= _GEN_4393;
      end
    end else begin
      data_9_0_4 <= _GEN_4393;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_5 <= _GEN_4457;
      end
    end else begin
      data_9_0_5 <= _GEN_4457;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_6 <= _GEN_4521;
      end
    end else begin
      data_9_0_6 <= _GEN_4521;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_0_7 <= _GEN_4585;
      end
    end else begin
      data_9_0_7 <= _GEN_4585;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_0 <= _GEN_4649;
      end
    end else begin
      data_9_1_0 <= _GEN_4649;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_1 <= _GEN_4713;
      end
    end else begin
      data_9_1_1 <= _GEN_4713;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_2 <= _GEN_4777;
      end
    end else begin
      data_9_1_2 <= _GEN_4777;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_3 <= _GEN_4841;
      end
    end else begin
      data_9_1_3 <= _GEN_4841;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_4 <= _GEN_4905;
      end
    end else begin
      data_9_1_4 <= _GEN_4905;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_5 <= _GEN_4969;
      end
    end else begin
      data_9_1_5 <= _GEN_4969;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_6 <= _GEN_5033;
      end
    end else begin
      data_9_1_6 <= _GEN_5033;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_1_7 <= _GEN_5097;
      end
    end else begin
      data_9_1_7 <= _GEN_5097;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_0 <= _GEN_5161;
      end
    end else begin
      data_9_2_0 <= _GEN_5161;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_1 <= _GEN_5225;
      end
    end else begin
      data_9_2_1 <= _GEN_5225;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_2 <= _GEN_5289;
      end
    end else begin
      data_9_2_2 <= _GEN_5289;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_3 <= _GEN_5353;
      end
    end else begin
      data_9_2_3 <= _GEN_5353;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_4 <= _GEN_5417;
      end
    end else begin
      data_9_2_4 <= _GEN_5417;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_5 <= _GEN_5481;
      end
    end else begin
      data_9_2_5 <= _GEN_5481;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_6 <= _GEN_5545;
      end
    end else begin
      data_9_2_6 <= _GEN_5545;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_2_7 <= _GEN_5609;
      end
    end else begin
      data_9_2_7 <= _GEN_5609;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_0 <= _GEN_5673;
      end
    end else begin
      data_9_3_0 <= _GEN_5673;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_1 <= _GEN_5737;
      end
    end else begin
      data_9_3_1 <= _GEN_5737;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_2 <= _GEN_5801;
      end
    end else begin
      data_9_3_2 <= _GEN_5801;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_3 <= _GEN_5865;
      end
    end else begin
      data_9_3_3 <= _GEN_5865;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_4 <= _GEN_5929;
      end
    end else begin
      data_9_3_4 <= _GEN_5929;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_5 <= _GEN_5993;
      end
    end else begin
      data_9_3_5 <= _GEN_5993;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_6 <= _GEN_6057;
      end
    end else begin
      data_9_3_6 <= _GEN_6057;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_3_7 <= _GEN_6121;
      end
    end else begin
      data_9_3_7 <= _GEN_6121;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_0 <= _GEN_6185;
      end
    end else begin
      data_9_4_0 <= _GEN_6185;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_1 <= _GEN_6249;
      end
    end else begin
      data_9_4_1 <= _GEN_6249;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_2 <= _GEN_6313;
      end
    end else begin
      data_9_4_2 <= _GEN_6313;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_3 <= _GEN_6377;
      end
    end else begin
      data_9_4_3 <= _GEN_6377;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_4 <= _GEN_6441;
      end
    end else begin
      data_9_4_4 <= _GEN_6441;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_5 <= _GEN_6505;
      end
    end else begin
      data_9_4_5 <= _GEN_6505;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_6 <= _GEN_6569;
      end
    end else begin
      data_9_4_6 <= _GEN_6569;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_4_7 <= _GEN_6633;
      end
    end else begin
      data_9_4_7 <= _GEN_6633;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_0 <= _GEN_6697;
      end
    end else begin
      data_9_5_0 <= _GEN_6697;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_1 <= _GEN_6761;
      end
    end else begin
      data_9_5_1 <= _GEN_6761;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_2 <= _GEN_6825;
      end
    end else begin
      data_9_5_2 <= _GEN_6825;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_3 <= _GEN_6889;
      end
    end else begin
      data_9_5_3 <= _GEN_6889;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_4 <= _GEN_6953;
      end
    end else begin
      data_9_5_4 <= _GEN_6953;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_5 <= _GEN_7017;
      end
    end else begin
      data_9_5_5 <= _GEN_7017;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_6 <= _GEN_7081;
      end
    end else begin
      data_9_5_6 <= _GEN_7081;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_5_7 <= _GEN_7145;
      end
    end else begin
      data_9_5_7 <= _GEN_7145;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_0 <= _GEN_7209;
      end
    end else begin
      data_9_6_0 <= _GEN_7209;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_1 <= _GEN_7273;
      end
    end else begin
      data_9_6_1 <= _GEN_7273;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_2 <= _GEN_7337;
      end
    end else begin
      data_9_6_2 <= _GEN_7337;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_3 <= _GEN_7401;
      end
    end else begin
      data_9_6_3 <= _GEN_7401;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_4 <= _GEN_7465;
      end
    end else begin
      data_9_6_4 <= _GEN_7465;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_5 <= _GEN_7529;
      end
    end else begin
      data_9_6_5 <= _GEN_7529;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_6 <= _GEN_7593;
      end
    end else begin
      data_9_6_6 <= _GEN_7593;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_6_7 <= _GEN_7657;
      end
    end else begin
      data_9_6_7 <= _GEN_7657;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_0 <= _GEN_7721;
      end
    end else begin
      data_9_7_0 <= _GEN_7721;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_1 <= _GEN_7785;
      end
    end else begin
      data_9_7_1 <= _GEN_7785;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_2 <= _GEN_7849;
      end
    end else begin
      data_9_7_2 <= _GEN_7849;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_3 <= _GEN_7913;
      end
    end else begin
      data_9_7_3 <= _GEN_7913;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_4 <= _GEN_7977;
      end
    end else begin
      data_9_7_4 <= _GEN_7977;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_5 <= _GEN_8041;
      end
    end else begin
      data_9_7_5 <= _GEN_8041;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_6 <= _GEN_8105;
      end
    end else begin
      data_9_7_6 <= _GEN_8105;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'h9 == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_9_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_9_7_7 <= _GEN_8169;
      end
    end else begin
      data_9_7_7 <= _GEN_8169;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_0 <= _GEN_4138;
      end
    end else begin
      data_10_0_0 <= _GEN_4138;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_1 <= _GEN_4202;
      end
    end else begin
      data_10_0_1 <= _GEN_4202;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_2 <= _GEN_4266;
      end
    end else begin
      data_10_0_2 <= _GEN_4266;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_3 <= _GEN_4330;
      end
    end else begin
      data_10_0_3 <= _GEN_4330;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_4 <= _GEN_4394;
      end
    end else begin
      data_10_0_4 <= _GEN_4394;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_5 <= _GEN_4458;
      end
    end else begin
      data_10_0_5 <= _GEN_4458;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_6 <= _GEN_4522;
      end
    end else begin
      data_10_0_6 <= _GEN_4522;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_0_7 <= _GEN_4586;
      end
    end else begin
      data_10_0_7 <= _GEN_4586;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_0 <= _GEN_4650;
      end
    end else begin
      data_10_1_0 <= _GEN_4650;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_1 <= _GEN_4714;
      end
    end else begin
      data_10_1_1 <= _GEN_4714;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_2 <= _GEN_4778;
      end
    end else begin
      data_10_1_2 <= _GEN_4778;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_3 <= _GEN_4842;
      end
    end else begin
      data_10_1_3 <= _GEN_4842;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_4 <= _GEN_4906;
      end
    end else begin
      data_10_1_4 <= _GEN_4906;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_5 <= _GEN_4970;
      end
    end else begin
      data_10_1_5 <= _GEN_4970;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_6 <= _GEN_5034;
      end
    end else begin
      data_10_1_6 <= _GEN_5034;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_1_7 <= _GEN_5098;
      end
    end else begin
      data_10_1_7 <= _GEN_5098;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_0 <= _GEN_5162;
      end
    end else begin
      data_10_2_0 <= _GEN_5162;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_1 <= _GEN_5226;
      end
    end else begin
      data_10_2_1 <= _GEN_5226;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_2 <= _GEN_5290;
      end
    end else begin
      data_10_2_2 <= _GEN_5290;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_3 <= _GEN_5354;
      end
    end else begin
      data_10_2_3 <= _GEN_5354;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_4 <= _GEN_5418;
      end
    end else begin
      data_10_2_4 <= _GEN_5418;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_5 <= _GEN_5482;
      end
    end else begin
      data_10_2_5 <= _GEN_5482;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_6 <= _GEN_5546;
      end
    end else begin
      data_10_2_6 <= _GEN_5546;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_2_7 <= _GEN_5610;
      end
    end else begin
      data_10_2_7 <= _GEN_5610;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_0 <= _GEN_5674;
      end
    end else begin
      data_10_3_0 <= _GEN_5674;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_1 <= _GEN_5738;
      end
    end else begin
      data_10_3_1 <= _GEN_5738;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_2 <= _GEN_5802;
      end
    end else begin
      data_10_3_2 <= _GEN_5802;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_3 <= _GEN_5866;
      end
    end else begin
      data_10_3_3 <= _GEN_5866;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_4 <= _GEN_5930;
      end
    end else begin
      data_10_3_4 <= _GEN_5930;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_5 <= _GEN_5994;
      end
    end else begin
      data_10_3_5 <= _GEN_5994;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_6 <= _GEN_6058;
      end
    end else begin
      data_10_3_6 <= _GEN_6058;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_3_7 <= _GEN_6122;
      end
    end else begin
      data_10_3_7 <= _GEN_6122;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_0 <= _GEN_6186;
      end
    end else begin
      data_10_4_0 <= _GEN_6186;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_1 <= _GEN_6250;
      end
    end else begin
      data_10_4_1 <= _GEN_6250;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_2 <= _GEN_6314;
      end
    end else begin
      data_10_4_2 <= _GEN_6314;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_3 <= _GEN_6378;
      end
    end else begin
      data_10_4_3 <= _GEN_6378;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_4 <= _GEN_6442;
      end
    end else begin
      data_10_4_4 <= _GEN_6442;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_5 <= _GEN_6506;
      end
    end else begin
      data_10_4_5 <= _GEN_6506;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_6 <= _GEN_6570;
      end
    end else begin
      data_10_4_6 <= _GEN_6570;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_4_7 <= _GEN_6634;
      end
    end else begin
      data_10_4_7 <= _GEN_6634;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_0 <= _GEN_6698;
      end
    end else begin
      data_10_5_0 <= _GEN_6698;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_1 <= _GEN_6762;
      end
    end else begin
      data_10_5_1 <= _GEN_6762;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_2 <= _GEN_6826;
      end
    end else begin
      data_10_5_2 <= _GEN_6826;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_3 <= _GEN_6890;
      end
    end else begin
      data_10_5_3 <= _GEN_6890;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_4 <= _GEN_6954;
      end
    end else begin
      data_10_5_4 <= _GEN_6954;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_5 <= _GEN_7018;
      end
    end else begin
      data_10_5_5 <= _GEN_7018;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_6 <= _GEN_7082;
      end
    end else begin
      data_10_5_6 <= _GEN_7082;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_5_7 <= _GEN_7146;
      end
    end else begin
      data_10_5_7 <= _GEN_7146;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_0 <= _GEN_7210;
      end
    end else begin
      data_10_6_0 <= _GEN_7210;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_1 <= _GEN_7274;
      end
    end else begin
      data_10_6_1 <= _GEN_7274;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_2 <= _GEN_7338;
      end
    end else begin
      data_10_6_2 <= _GEN_7338;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_3 <= _GEN_7402;
      end
    end else begin
      data_10_6_3 <= _GEN_7402;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_4 <= _GEN_7466;
      end
    end else begin
      data_10_6_4 <= _GEN_7466;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_5 <= _GEN_7530;
      end
    end else begin
      data_10_6_5 <= _GEN_7530;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_6 <= _GEN_7594;
      end
    end else begin
      data_10_6_6 <= _GEN_7594;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_6_7 <= _GEN_7658;
      end
    end else begin
      data_10_6_7 <= _GEN_7658;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_0 <= _GEN_7722;
      end
    end else begin
      data_10_7_0 <= _GEN_7722;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_1 <= _GEN_7786;
      end
    end else begin
      data_10_7_1 <= _GEN_7786;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_2 <= _GEN_7850;
      end
    end else begin
      data_10_7_2 <= _GEN_7850;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_3 <= _GEN_7914;
      end
    end else begin
      data_10_7_3 <= _GEN_7914;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_4 <= _GEN_7978;
      end
    end else begin
      data_10_7_4 <= _GEN_7978;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_5 <= _GEN_8042;
      end
    end else begin
      data_10_7_5 <= _GEN_8042;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_6 <= _GEN_8106;
      end
    end else begin
      data_10_7_6 <= _GEN_8106;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'ha == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_10_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_10_7_7 <= _GEN_8170;
      end
    end else begin
      data_10_7_7 <= _GEN_8170;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_0 <= _GEN_4139;
      end
    end else begin
      data_11_0_0 <= _GEN_4139;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_1 <= _GEN_4203;
      end
    end else begin
      data_11_0_1 <= _GEN_4203;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_2 <= _GEN_4267;
      end
    end else begin
      data_11_0_2 <= _GEN_4267;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_3 <= _GEN_4331;
      end
    end else begin
      data_11_0_3 <= _GEN_4331;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_4 <= _GEN_4395;
      end
    end else begin
      data_11_0_4 <= _GEN_4395;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_5 <= _GEN_4459;
      end
    end else begin
      data_11_0_5 <= _GEN_4459;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_6 <= _GEN_4523;
      end
    end else begin
      data_11_0_6 <= _GEN_4523;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_0_7 <= _GEN_4587;
      end
    end else begin
      data_11_0_7 <= _GEN_4587;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_0 <= _GEN_4651;
      end
    end else begin
      data_11_1_0 <= _GEN_4651;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_1 <= _GEN_4715;
      end
    end else begin
      data_11_1_1 <= _GEN_4715;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_2 <= _GEN_4779;
      end
    end else begin
      data_11_1_2 <= _GEN_4779;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_3 <= _GEN_4843;
      end
    end else begin
      data_11_1_3 <= _GEN_4843;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_4 <= _GEN_4907;
      end
    end else begin
      data_11_1_4 <= _GEN_4907;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_5 <= _GEN_4971;
      end
    end else begin
      data_11_1_5 <= _GEN_4971;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_6 <= _GEN_5035;
      end
    end else begin
      data_11_1_6 <= _GEN_5035;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_1_7 <= _GEN_5099;
      end
    end else begin
      data_11_1_7 <= _GEN_5099;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_0 <= _GEN_5163;
      end
    end else begin
      data_11_2_0 <= _GEN_5163;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_1 <= _GEN_5227;
      end
    end else begin
      data_11_2_1 <= _GEN_5227;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_2 <= _GEN_5291;
      end
    end else begin
      data_11_2_2 <= _GEN_5291;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_3 <= _GEN_5355;
      end
    end else begin
      data_11_2_3 <= _GEN_5355;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_4 <= _GEN_5419;
      end
    end else begin
      data_11_2_4 <= _GEN_5419;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_5 <= _GEN_5483;
      end
    end else begin
      data_11_2_5 <= _GEN_5483;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_6 <= _GEN_5547;
      end
    end else begin
      data_11_2_6 <= _GEN_5547;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_2_7 <= _GEN_5611;
      end
    end else begin
      data_11_2_7 <= _GEN_5611;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_0 <= _GEN_5675;
      end
    end else begin
      data_11_3_0 <= _GEN_5675;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_1 <= _GEN_5739;
      end
    end else begin
      data_11_3_1 <= _GEN_5739;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_2 <= _GEN_5803;
      end
    end else begin
      data_11_3_2 <= _GEN_5803;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_3 <= _GEN_5867;
      end
    end else begin
      data_11_3_3 <= _GEN_5867;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_4 <= _GEN_5931;
      end
    end else begin
      data_11_3_4 <= _GEN_5931;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_5 <= _GEN_5995;
      end
    end else begin
      data_11_3_5 <= _GEN_5995;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_6 <= _GEN_6059;
      end
    end else begin
      data_11_3_6 <= _GEN_6059;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_3_7 <= _GEN_6123;
      end
    end else begin
      data_11_3_7 <= _GEN_6123;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_0 <= _GEN_6187;
      end
    end else begin
      data_11_4_0 <= _GEN_6187;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_1 <= _GEN_6251;
      end
    end else begin
      data_11_4_1 <= _GEN_6251;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_2 <= _GEN_6315;
      end
    end else begin
      data_11_4_2 <= _GEN_6315;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_3 <= _GEN_6379;
      end
    end else begin
      data_11_4_3 <= _GEN_6379;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_4 <= _GEN_6443;
      end
    end else begin
      data_11_4_4 <= _GEN_6443;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_5 <= _GEN_6507;
      end
    end else begin
      data_11_4_5 <= _GEN_6507;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_6 <= _GEN_6571;
      end
    end else begin
      data_11_4_6 <= _GEN_6571;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_4_7 <= _GEN_6635;
      end
    end else begin
      data_11_4_7 <= _GEN_6635;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_0 <= _GEN_6699;
      end
    end else begin
      data_11_5_0 <= _GEN_6699;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_1 <= _GEN_6763;
      end
    end else begin
      data_11_5_1 <= _GEN_6763;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_2 <= _GEN_6827;
      end
    end else begin
      data_11_5_2 <= _GEN_6827;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_3 <= _GEN_6891;
      end
    end else begin
      data_11_5_3 <= _GEN_6891;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_4 <= _GEN_6955;
      end
    end else begin
      data_11_5_4 <= _GEN_6955;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_5 <= _GEN_7019;
      end
    end else begin
      data_11_5_5 <= _GEN_7019;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_6 <= _GEN_7083;
      end
    end else begin
      data_11_5_6 <= _GEN_7083;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_5_7 <= _GEN_7147;
      end
    end else begin
      data_11_5_7 <= _GEN_7147;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_0 <= _GEN_7211;
      end
    end else begin
      data_11_6_0 <= _GEN_7211;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_1 <= _GEN_7275;
      end
    end else begin
      data_11_6_1 <= _GEN_7275;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_2 <= _GEN_7339;
      end
    end else begin
      data_11_6_2 <= _GEN_7339;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_3 <= _GEN_7403;
      end
    end else begin
      data_11_6_3 <= _GEN_7403;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_4 <= _GEN_7467;
      end
    end else begin
      data_11_6_4 <= _GEN_7467;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_5 <= _GEN_7531;
      end
    end else begin
      data_11_6_5 <= _GEN_7531;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_6 <= _GEN_7595;
      end
    end else begin
      data_11_6_6 <= _GEN_7595;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_6_7 <= _GEN_7659;
      end
    end else begin
      data_11_6_7 <= _GEN_7659;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_0 <= _GEN_7723;
      end
    end else begin
      data_11_7_0 <= _GEN_7723;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_1 <= _GEN_7787;
      end
    end else begin
      data_11_7_1 <= _GEN_7787;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_2 <= _GEN_7851;
      end
    end else begin
      data_11_7_2 <= _GEN_7851;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_3 <= _GEN_7915;
      end
    end else begin
      data_11_7_3 <= _GEN_7915;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_4 <= _GEN_7979;
      end
    end else begin
      data_11_7_4 <= _GEN_7979;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_5 <= _GEN_8043;
      end
    end else begin
      data_11_7_5 <= _GEN_8043;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_6 <= _GEN_8107;
      end
    end else begin
      data_11_7_6 <= _GEN_8107;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'hb == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_11_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_11_7_7 <= _GEN_8171;
      end
    end else begin
      data_11_7_7 <= _GEN_8171;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_0 <= _GEN_4140;
      end
    end else begin
      data_12_0_0 <= _GEN_4140;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_1 <= _GEN_4204;
      end
    end else begin
      data_12_0_1 <= _GEN_4204;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_2 <= _GEN_4268;
      end
    end else begin
      data_12_0_2 <= _GEN_4268;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_3 <= _GEN_4332;
      end
    end else begin
      data_12_0_3 <= _GEN_4332;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_4 <= _GEN_4396;
      end
    end else begin
      data_12_0_4 <= _GEN_4396;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_5 <= _GEN_4460;
      end
    end else begin
      data_12_0_5 <= _GEN_4460;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_6 <= _GEN_4524;
      end
    end else begin
      data_12_0_6 <= _GEN_4524;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_0_7 <= _GEN_4588;
      end
    end else begin
      data_12_0_7 <= _GEN_4588;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_0 <= _GEN_4652;
      end
    end else begin
      data_12_1_0 <= _GEN_4652;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_1 <= _GEN_4716;
      end
    end else begin
      data_12_1_1 <= _GEN_4716;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_2 <= _GEN_4780;
      end
    end else begin
      data_12_1_2 <= _GEN_4780;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_3 <= _GEN_4844;
      end
    end else begin
      data_12_1_3 <= _GEN_4844;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_4 <= _GEN_4908;
      end
    end else begin
      data_12_1_4 <= _GEN_4908;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_5 <= _GEN_4972;
      end
    end else begin
      data_12_1_5 <= _GEN_4972;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_6 <= _GEN_5036;
      end
    end else begin
      data_12_1_6 <= _GEN_5036;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_1_7 <= _GEN_5100;
      end
    end else begin
      data_12_1_7 <= _GEN_5100;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_0 <= _GEN_5164;
      end
    end else begin
      data_12_2_0 <= _GEN_5164;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_1 <= _GEN_5228;
      end
    end else begin
      data_12_2_1 <= _GEN_5228;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_2 <= _GEN_5292;
      end
    end else begin
      data_12_2_2 <= _GEN_5292;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_3 <= _GEN_5356;
      end
    end else begin
      data_12_2_3 <= _GEN_5356;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_4 <= _GEN_5420;
      end
    end else begin
      data_12_2_4 <= _GEN_5420;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_5 <= _GEN_5484;
      end
    end else begin
      data_12_2_5 <= _GEN_5484;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_6 <= _GEN_5548;
      end
    end else begin
      data_12_2_6 <= _GEN_5548;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_2_7 <= _GEN_5612;
      end
    end else begin
      data_12_2_7 <= _GEN_5612;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_0 <= _GEN_5676;
      end
    end else begin
      data_12_3_0 <= _GEN_5676;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_1 <= _GEN_5740;
      end
    end else begin
      data_12_3_1 <= _GEN_5740;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_2 <= _GEN_5804;
      end
    end else begin
      data_12_3_2 <= _GEN_5804;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_3 <= _GEN_5868;
      end
    end else begin
      data_12_3_3 <= _GEN_5868;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_4 <= _GEN_5932;
      end
    end else begin
      data_12_3_4 <= _GEN_5932;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_5 <= _GEN_5996;
      end
    end else begin
      data_12_3_5 <= _GEN_5996;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_6 <= _GEN_6060;
      end
    end else begin
      data_12_3_6 <= _GEN_6060;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_3_7 <= _GEN_6124;
      end
    end else begin
      data_12_3_7 <= _GEN_6124;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_0 <= _GEN_6188;
      end
    end else begin
      data_12_4_0 <= _GEN_6188;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_1 <= _GEN_6252;
      end
    end else begin
      data_12_4_1 <= _GEN_6252;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_2 <= _GEN_6316;
      end
    end else begin
      data_12_4_2 <= _GEN_6316;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_3 <= _GEN_6380;
      end
    end else begin
      data_12_4_3 <= _GEN_6380;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_4 <= _GEN_6444;
      end
    end else begin
      data_12_4_4 <= _GEN_6444;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_5 <= _GEN_6508;
      end
    end else begin
      data_12_4_5 <= _GEN_6508;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_6 <= _GEN_6572;
      end
    end else begin
      data_12_4_6 <= _GEN_6572;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_4_7 <= _GEN_6636;
      end
    end else begin
      data_12_4_7 <= _GEN_6636;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_0 <= _GEN_6700;
      end
    end else begin
      data_12_5_0 <= _GEN_6700;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_1 <= _GEN_6764;
      end
    end else begin
      data_12_5_1 <= _GEN_6764;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_2 <= _GEN_6828;
      end
    end else begin
      data_12_5_2 <= _GEN_6828;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_3 <= _GEN_6892;
      end
    end else begin
      data_12_5_3 <= _GEN_6892;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_4 <= _GEN_6956;
      end
    end else begin
      data_12_5_4 <= _GEN_6956;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_5 <= _GEN_7020;
      end
    end else begin
      data_12_5_5 <= _GEN_7020;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_6 <= _GEN_7084;
      end
    end else begin
      data_12_5_6 <= _GEN_7084;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_5_7 <= _GEN_7148;
      end
    end else begin
      data_12_5_7 <= _GEN_7148;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_0 <= _GEN_7212;
      end
    end else begin
      data_12_6_0 <= _GEN_7212;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_1 <= _GEN_7276;
      end
    end else begin
      data_12_6_1 <= _GEN_7276;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_2 <= _GEN_7340;
      end
    end else begin
      data_12_6_2 <= _GEN_7340;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_3 <= _GEN_7404;
      end
    end else begin
      data_12_6_3 <= _GEN_7404;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_4 <= _GEN_7468;
      end
    end else begin
      data_12_6_4 <= _GEN_7468;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_5 <= _GEN_7532;
      end
    end else begin
      data_12_6_5 <= _GEN_7532;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_6 <= _GEN_7596;
      end
    end else begin
      data_12_6_6 <= _GEN_7596;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_6_7 <= _GEN_7660;
      end
    end else begin
      data_12_6_7 <= _GEN_7660;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_0 <= _GEN_7724;
      end
    end else begin
      data_12_7_0 <= _GEN_7724;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_1 <= _GEN_7788;
      end
    end else begin
      data_12_7_1 <= _GEN_7788;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_2 <= _GEN_7852;
      end
    end else begin
      data_12_7_2 <= _GEN_7852;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_3 <= _GEN_7916;
      end
    end else begin
      data_12_7_3 <= _GEN_7916;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_4 <= _GEN_7980;
      end
    end else begin
      data_12_7_4 <= _GEN_7980;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_5 <= _GEN_8044;
      end
    end else begin
      data_12_7_5 <= _GEN_8044;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_6 <= _GEN_8108;
      end
    end else begin
      data_12_7_6 <= _GEN_8108;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'hc == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_12_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_12_7_7 <= _GEN_8172;
      end
    end else begin
      data_12_7_7 <= _GEN_8172;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_0 <= _GEN_4141;
      end
    end else begin
      data_13_0_0 <= _GEN_4141;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_1 <= _GEN_4205;
      end
    end else begin
      data_13_0_1 <= _GEN_4205;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_2 <= _GEN_4269;
      end
    end else begin
      data_13_0_2 <= _GEN_4269;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_3 <= _GEN_4333;
      end
    end else begin
      data_13_0_3 <= _GEN_4333;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_4 <= _GEN_4397;
      end
    end else begin
      data_13_0_4 <= _GEN_4397;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_5 <= _GEN_4461;
      end
    end else begin
      data_13_0_5 <= _GEN_4461;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_6 <= _GEN_4525;
      end
    end else begin
      data_13_0_6 <= _GEN_4525;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_0_7 <= _GEN_4589;
      end
    end else begin
      data_13_0_7 <= _GEN_4589;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_0 <= _GEN_4653;
      end
    end else begin
      data_13_1_0 <= _GEN_4653;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_1 <= _GEN_4717;
      end
    end else begin
      data_13_1_1 <= _GEN_4717;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_2 <= _GEN_4781;
      end
    end else begin
      data_13_1_2 <= _GEN_4781;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_3 <= _GEN_4845;
      end
    end else begin
      data_13_1_3 <= _GEN_4845;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_4 <= _GEN_4909;
      end
    end else begin
      data_13_1_4 <= _GEN_4909;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_5 <= _GEN_4973;
      end
    end else begin
      data_13_1_5 <= _GEN_4973;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_6 <= _GEN_5037;
      end
    end else begin
      data_13_1_6 <= _GEN_5037;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_1_7 <= _GEN_5101;
      end
    end else begin
      data_13_1_7 <= _GEN_5101;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_0 <= _GEN_5165;
      end
    end else begin
      data_13_2_0 <= _GEN_5165;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_1 <= _GEN_5229;
      end
    end else begin
      data_13_2_1 <= _GEN_5229;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_2 <= _GEN_5293;
      end
    end else begin
      data_13_2_2 <= _GEN_5293;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_3 <= _GEN_5357;
      end
    end else begin
      data_13_2_3 <= _GEN_5357;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_4 <= _GEN_5421;
      end
    end else begin
      data_13_2_4 <= _GEN_5421;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_5 <= _GEN_5485;
      end
    end else begin
      data_13_2_5 <= _GEN_5485;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_6 <= _GEN_5549;
      end
    end else begin
      data_13_2_6 <= _GEN_5549;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_2_7 <= _GEN_5613;
      end
    end else begin
      data_13_2_7 <= _GEN_5613;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_0 <= _GEN_5677;
      end
    end else begin
      data_13_3_0 <= _GEN_5677;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_1 <= _GEN_5741;
      end
    end else begin
      data_13_3_1 <= _GEN_5741;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_2 <= _GEN_5805;
      end
    end else begin
      data_13_3_2 <= _GEN_5805;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_3 <= _GEN_5869;
      end
    end else begin
      data_13_3_3 <= _GEN_5869;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_4 <= _GEN_5933;
      end
    end else begin
      data_13_3_4 <= _GEN_5933;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_5 <= _GEN_5997;
      end
    end else begin
      data_13_3_5 <= _GEN_5997;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_6 <= _GEN_6061;
      end
    end else begin
      data_13_3_6 <= _GEN_6061;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_3_7 <= _GEN_6125;
      end
    end else begin
      data_13_3_7 <= _GEN_6125;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_0 <= _GEN_6189;
      end
    end else begin
      data_13_4_0 <= _GEN_6189;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_1 <= _GEN_6253;
      end
    end else begin
      data_13_4_1 <= _GEN_6253;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_2 <= _GEN_6317;
      end
    end else begin
      data_13_4_2 <= _GEN_6317;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_3 <= _GEN_6381;
      end
    end else begin
      data_13_4_3 <= _GEN_6381;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_4 <= _GEN_6445;
      end
    end else begin
      data_13_4_4 <= _GEN_6445;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_5 <= _GEN_6509;
      end
    end else begin
      data_13_4_5 <= _GEN_6509;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_6 <= _GEN_6573;
      end
    end else begin
      data_13_4_6 <= _GEN_6573;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_4_7 <= _GEN_6637;
      end
    end else begin
      data_13_4_7 <= _GEN_6637;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_0 <= _GEN_6701;
      end
    end else begin
      data_13_5_0 <= _GEN_6701;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_1 <= _GEN_6765;
      end
    end else begin
      data_13_5_1 <= _GEN_6765;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_2 <= _GEN_6829;
      end
    end else begin
      data_13_5_2 <= _GEN_6829;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_3 <= _GEN_6893;
      end
    end else begin
      data_13_5_3 <= _GEN_6893;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_4 <= _GEN_6957;
      end
    end else begin
      data_13_5_4 <= _GEN_6957;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_5 <= _GEN_7021;
      end
    end else begin
      data_13_5_5 <= _GEN_7021;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_6 <= _GEN_7085;
      end
    end else begin
      data_13_5_6 <= _GEN_7085;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_5_7 <= _GEN_7149;
      end
    end else begin
      data_13_5_7 <= _GEN_7149;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_0 <= _GEN_7213;
      end
    end else begin
      data_13_6_0 <= _GEN_7213;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_1 <= _GEN_7277;
      end
    end else begin
      data_13_6_1 <= _GEN_7277;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_2 <= _GEN_7341;
      end
    end else begin
      data_13_6_2 <= _GEN_7341;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_3 <= _GEN_7405;
      end
    end else begin
      data_13_6_3 <= _GEN_7405;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_4 <= _GEN_7469;
      end
    end else begin
      data_13_6_4 <= _GEN_7469;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_5 <= _GEN_7533;
      end
    end else begin
      data_13_6_5 <= _GEN_7533;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_6 <= _GEN_7597;
      end
    end else begin
      data_13_6_6 <= _GEN_7597;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_6_7 <= _GEN_7661;
      end
    end else begin
      data_13_6_7 <= _GEN_7661;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_0 <= _GEN_7725;
      end
    end else begin
      data_13_7_0 <= _GEN_7725;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_1 <= _GEN_7789;
      end
    end else begin
      data_13_7_1 <= _GEN_7789;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_2 <= _GEN_7853;
      end
    end else begin
      data_13_7_2 <= _GEN_7853;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_3 <= _GEN_7917;
      end
    end else begin
      data_13_7_3 <= _GEN_7917;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_4 <= _GEN_7981;
      end
    end else begin
      data_13_7_4 <= _GEN_7981;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_5 <= _GEN_8045;
      end
    end else begin
      data_13_7_5 <= _GEN_8045;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_6 <= _GEN_8109;
      end
    end else begin
      data_13_7_6 <= _GEN_8109;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'hd == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_13_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_13_7_7 <= _GEN_8173;
      end
    end else begin
      data_13_7_7 <= _GEN_8173;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_0 <= _GEN_4142;
      end
    end else begin
      data_14_0_0 <= _GEN_4142;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_1 <= _GEN_4206;
      end
    end else begin
      data_14_0_1 <= _GEN_4206;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_2 <= _GEN_4270;
      end
    end else begin
      data_14_0_2 <= _GEN_4270;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_3 <= _GEN_4334;
      end
    end else begin
      data_14_0_3 <= _GEN_4334;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_4 <= _GEN_4398;
      end
    end else begin
      data_14_0_4 <= _GEN_4398;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_5 <= _GEN_4462;
      end
    end else begin
      data_14_0_5 <= _GEN_4462;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_6 <= _GEN_4526;
      end
    end else begin
      data_14_0_6 <= _GEN_4526;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_0_7 <= _GEN_4590;
      end
    end else begin
      data_14_0_7 <= _GEN_4590;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_0 <= _GEN_4654;
      end
    end else begin
      data_14_1_0 <= _GEN_4654;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_1 <= _GEN_4718;
      end
    end else begin
      data_14_1_1 <= _GEN_4718;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_2 <= _GEN_4782;
      end
    end else begin
      data_14_1_2 <= _GEN_4782;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_3 <= _GEN_4846;
      end
    end else begin
      data_14_1_3 <= _GEN_4846;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_4 <= _GEN_4910;
      end
    end else begin
      data_14_1_4 <= _GEN_4910;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_5 <= _GEN_4974;
      end
    end else begin
      data_14_1_5 <= _GEN_4974;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_6 <= _GEN_5038;
      end
    end else begin
      data_14_1_6 <= _GEN_5038;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_1_7 <= _GEN_5102;
      end
    end else begin
      data_14_1_7 <= _GEN_5102;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_0 <= _GEN_5166;
      end
    end else begin
      data_14_2_0 <= _GEN_5166;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_1 <= _GEN_5230;
      end
    end else begin
      data_14_2_1 <= _GEN_5230;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_2 <= _GEN_5294;
      end
    end else begin
      data_14_2_2 <= _GEN_5294;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_3 <= _GEN_5358;
      end
    end else begin
      data_14_2_3 <= _GEN_5358;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_4 <= _GEN_5422;
      end
    end else begin
      data_14_2_4 <= _GEN_5422;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_5 <= _GEN_5486;
      end
    end else begin
      data_14_2_5 <= _GEN_5486;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_6 <= _GEN_5550;
      end
    end else begin
      data_14_2_6 <= _GEN_5550;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_2_7 <= _GEN_5614;
      end
    end else begin
      data_14_2_7 <= _GEN_5614;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_0 <= _GEN_5678;
      end
    end else begin
      data_14_3_0 <= _GEN_5678;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_1 <= _GEN_5742;
      end
    end else begin
      data_14_3_1 <= _GEN_5742;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_2 <= _GEN_5806;
      end
    end else begin
      data_14_3_2 <= _GEN_5806;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_3 <= _GEN_5870;
      end
    end else begin
      data_14_3_3 <= _GEN_5870;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_4 <= _GEN_5934;
      end
    end else begin
      data_14_3_4 <= _GEN_5934;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_5 <= _GEN_5998;
      end
    end else begin
      data_14_3_5 <= _GEN_5998;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_6 <= _GEN_6062;
      end
    end else begin
      data_14_3_6 <= _GEN_6062;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_3_7 <= _GEN_6126;
      end
    end else begin
      data_14_3_7 <= _GEN_6126;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_0 <= _GEN_6190;
      end
    end else begin
      data_14_4_0 <= _GEN_6190;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_1 <= _GEN_6254;
      end
    end else begin
      data_14_4_1 <= _GEN_6254;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_2 <= _GEN_6318;
      end
    end else begin
      data_14_4_2 <= _GEN_6318;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_3 <= _GEN_6382;
      end
    end else begin
      data_14_4_3 <= _GEN_6382;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_4 <= _GEN_6446;
      end
    end else begin
      data_14_4_4 <= _GEN_6446;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_5 <= _GEN_6510;
      end
    end else begin
      data_14_4_5 <= _GEN_6510;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_6 <= _GEN_6574;
      end
    end else begin
      data_14_4_6 <= _GEN_6574;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_4_7 <= _GEN_6638;
      end
    end else begin
      data_14_4_7 <= _GEN_6638;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_0 <= _GEN_6702;
      end
    end else begin
      data_14_5_0 <= _GEN_6702;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_1 <= _GEN_6766;
      end
    end else begin
      data_14_5_1 <= _GEN_6766;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_2 <= _GEN_6830;
      end
    end else begin
      data_14_5_2 <= _GEN_6830;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_3 <= _GEN_6894;
      end
    end else begin
      data_14_5_3 <= _GEN_6894;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_4 <= _GEN_6958;
      end
    end else begin
      data_14_5_4 <= _GEN_6958;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_5 <= _GEN_7022;
      end
    end else begin
      data_14_5_5 <= _GEN_7022;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_6 <= _GEN_7086;
      end
    end else begin
      data_14_5_6 <= _GEN_7086;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_5_7 <= _GEN_7150;
      end
    end else begin
      data_14_5_7 <= _GEN_7150;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_0 <= _GEN_7214;
      end
    end else begin
      data_14_6_0 <= _GEN_7214;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_1 <= _GEN_7278;
      end
    end else begin
      data_14_6_1 <= _GEN_7278;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_2 <= _GEN_7342;
      end
    end else begin
      data_14_6_2 <= _GEN_7342;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_3 <= _GEN_7406;
      end
    end else begin
      data_14_6_3 <= _GEN_7406;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_4 <= _GEN_7470;
      end
    end else begin
      data_14_6_4 <= _GEN_7470;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_5 <= _GEN_7534;
      end
    end else begin
      data_14_6_5 <= _GEN_7534;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_6 <= _GEN_7598;
      end
    end else begin
      data_14_6_6 <= _GEN_7598;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_6_7 <= _GEN_7662;
      end
    end else begin
      data_14_6_7 <= _GEN_7662;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_0 <= _GEN_7726;
      end
    end else begin
      data_14_7_0 <= _GEN_7726;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_1 <= _GEN_7790;
      end
    end else begin
      data_14_7_1 <= _GEN_7790;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_2 <= _GEN_7854;
      end
    end else begin
      data_14_7_2 <= _GEN_7854;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_3 <= _GEN_7918;
      end
    end else begin
      data_14_7_3 <= _GEN_7918;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_4 <= _GEN_7982;
      end
    end else begin
      data_14_7_4 <= _GEN_7982;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_5 <= _GEN_8046;
      end
    end else begin
      data_14_7_5 <= _GEN_8046;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_6 <= _GEN_8110;
      end
    end else begin
      data_14_7_6 <= _GEN_8110;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'he == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_14_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_14_7_7 <= _GEN_8174;
      end
    end else begin
      data_14_7_7 <= _GEN_8174;
    end
    if (wen_64) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_0 <= _GEN_4143;
      end
    end else begin
      data_15_0_0 <= _GEN_4143;
    end
    if (wen_65) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_1 <= _GEN_4207;
      end
    end else begin
      data_15_0_1 <= _GEN_4207;
    end
    if (wen_66) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_2 <= _GEN_4271;
      end
    end else begin
      data_15_0_2 <= _GEN_4271;
    end
    if (wen_67) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_3 <= _GEN_4335;
      end
    end else begin
      data_15_0_3 <= _GEN_4335;
    end
    if (wen_68) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_4 <= _GEN_4399;
      end
    end else begin
      data_15_0_4 <= _GEN_4399;
    end
    if (wen_69) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_5 <= _GEN_4463;
      end
    end else begin
      data_15_0_5 <= _GEN_4463;
    end
    if (wen_70) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_6 <= _GEN_4527;
      end
    end else begin
      data_15_0_6 <= _GEN_4527;
    end
    if (wen_71) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_0_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_0_7 <= _GEN_4591;
      end
    end else begin
      data_15_0_7 <= _GEN_4591;
    end
    if (wen_72) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_0 <= _GEN_4655;
      end
    end else begin
      data_15_1_0 <= _GEN_4655;
    end
    if (wen_73) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_1 <= _GEN_4719;
      end
    end else begin
      data_15_1_1 <= _GEN_4719;
    end
    if (wen_74) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_2 <= _GEN_4783;
      end
    end else begin
      data_15_1_2 <= _GEN_4783;
    end
    if (wen_75) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_3 <= _GEN_4847;
      end
    end else begin
      data_15_1_3 <= _GEN_4847;
    end
    if (wen_76) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_4 <= _GEN_4911;
      end
    end else begin
      data_15_1_4 <= _GEN_4911;
    end
    if (wen_77) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_5 <= _GEN_4975;
      end
    end else begin
      data_15_1_5 <= _GEN_4975;
    end
    if (wen_78) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_6 <= _GEN_5039;
      end
    end else begin
      data_15_1_6 <= _GEN_5039;
    end
    if (wen_79) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_1_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_1_7 <= _GEN_5103;
      end
    end else begin
      data_15_1_7 <= _GEN_5103;
    end
    if (wen_80) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_0 <= _GEN_5167;
      end
    end else begin
      data_15_2_0 <= _GEN_5167;
    end
    if (wen_81) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_1 <= _GEN_5231;
      end
    end else begin
      data_15_2_1 <= _GEN_5231;
    end
    if (wen_82) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_2 <= _GEN_5295;
      end
    end else begin
      data_15_2_2 <= _GEN_5295;
    end
    if (wen_83) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_3 <= _GEN_5359;
      end
    end else begin
      data_15_2_3 <= _GEN_5359;
    end
    if (wen_84) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_4 <= _GEN_5423;
      end
    end else begin
      data_15_2_4 <= _GEN_5423;
    end
    if (wen_85) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_5 <= _GEN_5487;
      end
    end else begin
      data_15_2_5 <= _GEN_5487;
    end
    if (wen_86) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_6 <= _GEN_5551;
      end
    end else begin
      data_15_2_6 <= _GEN_5551;
    end
    if (wen_87) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_2_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_2_7 <= _GEN_5615;
      end
    end else begin
      data_15_2_7 <= _GEN_5615;
    end
    if (wen_88) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_0 <= _GEN_5679;
      end
    end else begin
      data_15_3_0 <= _GEN_5679;
    end
    if (wen_89) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_1 <= _GEN_5743;
      end
    end else begin
      data_15_3_1 <= _GEN_5743;
    end
    if (wen_90) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_2 <= _GEN_5807;
      end
    end else begin
      data_15_3_2 <= _GEN_5807;
    end
    if (wen_91) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_3 <= _GEN_5871;
      end
    end else begin
      data_15_3_3 <= _GEN_5871;
    end
    if (wen_92) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_4 <= _GEN_5935;
      end
    end else begin
      data_15_3_4 <= _GEN_5935;
    end
    if (wen_93) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_5 <= _GEN_5999;
      end
    end else begin
      data_15_3_5 <= _GEN_5999;
    end
    if (wen_94) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_6 <= _GEN_6063;
      end
    end else begin
      data_15_3_6 <= _GEN_6063;
    end
    if (wen_95) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_3_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_3_7 <= _GEN_6127;
      end
    end else begin
      data_15_3_7 <= _GEN_6127;
    end
    if (wen_96) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_0 <= _GEN_6191;
      end
    end else begin
      data_15_4_0 <= _GEN_6191;
    end
    if (wen_97) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_1 <= _GEN_6255;
      end
    end else begin
      data_15_4_1 <= _GEN_6255;
    end
    if (wen_98) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_2 <= _GEN_6319;
      end
    end else begin
      data_15_4_2 <= _GEN_6319;
    end
    if (wen_99) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_3 <= _GEN_6383;
      end
    end else begin
      data_15_4_3 <= _GEN_6383;
    end
    if (wen_100) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_4 <= _GEN_6447;
      end
    end else begin
      data_15_4_4 <= _GEN_6447;
    end
    if (wen_101) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_5 <= _GEN_6511;
      end
    end else begin
      data_15_4_5 <= _GEN_6511;
    end
    if (wen_102) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_6 <= _GEN_6575;
      end
    end else begin
      data_15_4_6 <= _GEN_6575;
    end
    if (wen_103) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_4_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_4_7 <= _GEN_6639;
      end
    end else begin
      data_15_4_7 <= _GEN_6639;
    end
    if (wen_104) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_0 <= _GEN_6703;
      end
    end else begin
      data_15_5_0 <= _GEN_6703;
    end
    if (wen_105) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_1 <= _GEN_6767;
      end
    end else begin
      data_15_5_1 <= _GEN_6767;
    end
    if (wen_106) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_2 <= _GEN_6831;
      end
    end else begin
      data_15_5_2 <= _GEN_6831;
    end
    if (wen_107) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_3 <= _GEN_6895;
      end
    end else begin
      data_15_5_3 <= _GEN_6895;
    end
    if (wen_108) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_4 <= _GEN_6959;
      end
    end else begin
      data_15_5_4 <= _GEN_6959;
    end
    if (wen_109) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_5 <= _GEN_7023;
      end
    end else begin
      data_15_5_5 <= _GEN_7023;
    end
    if (wen_110) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_6 <= _GEN_7087;
      end
    end else begin
      data_15_5_6 <= _GEN_7087;
    end
    if (wen_111) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_5_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_5_7 <= _GEN_7151;
      end
    end else begin
      data_15_5_7 <= _GEN_7151;
    end
    if (wen_112) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_0 <= _GEN_7215;
      end
    end else begin
      data_15_6_0 <= _GEN_7215;
    end
    if (wen_113) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_1 <= _GEN_7279;
      end
    end else begin
      data_15_6_1 <= _GEN_7279;
    end
    if (wen_114) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_2 <= _GEN_7343;
      end
    end else begin
      data_15_6_2 <= _GEN_7343;
    end
    if (wen_115) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_3 <= _GEN_7407;
      end
    end else begin
      data_15_6_3 <= _GEN_7407;
    end
    if (wen_116) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_4 <= _GEN_7471;
      end
    end else begin
      data_15_6_4 <= _GEN_7471;
    end
    if (wen_117) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_5 <= _GEN_7535;
      end
    end else begin
      data_15_6_5 <= _GEN_7535;
    end
    if (wen_118) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_6 <= _GEN_7599;
      end
    end else begin
      data_15_6_6 <= _GEN_7599;
    end
    if (wen_119) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_6_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_6_7 <= _GEN_7663;
      end
    end else begin
      data_15_6_7 <= _GEN_7663;
    end
    if (wen_120) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_0 <= w_data_s1_1[7:0]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_0 <= _GEN_7727;
      end
    end else begin
      data_15_7_0 <= _GEN_7727;
    end
    if (wen_121) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_1 <= w_data_s1_1[15:8]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_1 <= _GEN_7791;
      end
    end else begin
      data_15_7_1 <= _GEN_7791;
    end
    if (wen_122) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_2 <= w_data_s1_1[23:16]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_2 <= _GEN_7855;
      end
    end else begin
      data_15_7_2 <= _GEN_7855;
    end
    if (wen_123) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_3 <= w_data_s1_1[31:24]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_3 <= _GEN_7919;
      end
    end else begin
      data_15_7_3 <= _GEN_7919;
    end
    if (wen_124) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_4 <= w_data_s1_1[39:32]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_4 <= _GEN_7983;
      end
    end else begin
      data_15_7_4 <= _GEN_7983;
    end
    if (wen_125) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_5 <= w_data_s1_1[47:40]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_5 <= _GEN_8047;
      end
    end else begin
      data_15_7_5 <= _GEN_8047;
    end
    if (wen_126) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_6 <= w_data_s1_1[55:48]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_6 <= _GEN_8111;
      end
    end else begin
      data_15_7_6 <= _GEN_8111;
    end
    if (wen_127) begin // @[Sbuffer.scala 160:18]
      if (4'hf == w_addr_s1_1) begin // @[Sbuffer.scala 161:42]
        data_15_7_7 <= w_data_s1_1[63:56]; // @[Sbuffer.scala 161:42]
      end else begin
        data_15_7_7 <= _GEN_8175;
      end
    end else begin
      data_15_7_7 <= _GEN_8175;
    end
    line_mask_clean_valid_0 <= io_maskFlushReq_0_valid; // @[Sbuffer.scala 121:63]
    line_mask_clean_valid_1 <= io_maskFlushReq_1_valid; // @[Sbuffer.scala 121:63]
    line_mask_clean_line_0 <= {_line_mask_clean_line_T,_line_mask_clean_line_T_8}; // @[Cat.scala 33:92]
    line_mask_clean_line_1 <= {_line_mask_clean_line_T_10,_line_mask_clean_line_T_18}; // @[Cat.scala 33:92]
    w_valid_s1_0 <= io_writeReq_0_valid; // @[Sbuffer.scala 146:40]
    w_valid_s1_1 <= io_writeReq_1_valid; // @[Sbuffer.scala 146:40]
    w_data_s1_0 <= io_writeReq_0_bits_data; // @[Sbuffer.scala 147:39]
    w_data_s1_1 <= io_writeReq_1_bits_data; // @[Sbuffer.scala 147:39]
    w_wline_s1_0 <= io_writeReq_0_bits_wline; // @[Sbuffer.scala 148:40]
    w_wline_s1_1 <= io_writeReq_1_bits_wline; // @[Sbuffer.scala 148:40]
    w_mask_s1_0 <= io_writeReq_0_bits_mask; // @[Sbuffer.scala 149:39]
    w_mask_s1_1 <= io_writeReq_1_bits_mask; // @[Sbuffer.scala 149:39]
    w_addr_s1_0 <= {_w_addr_s1_T,_w_addr_s1_T_8}; // @[Cat.scala 33:92]
    w_addr_s1_1 <= {_w_addr_s1_T_10,_w_addr_s1_T_18}; // @[Cat.scala 33:92]
    w_word_offset_s1_0 <= io_writeReq_0_bits_wordOffset[2:0]; // @[Sbuffer.scala 151:64]
    w_word_offset_s1_1 <= io_writeReq_1_bits_wordOffset[2:0]; // @[Sbuffer.scala 151:64]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_0_0_0 <= _GEN_8208;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_0_0_0 <= _GEN_4112; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_0 <= 1'h0;
      end else begin
        mask_0_0_0 <= _GEN_1024;
      end
    end else begin
      mask_0_0_0 <= _GEN_1024;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_0_0_1 <= _GEN_8272;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_0_0_1 <= _GEN_4176; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_1 <= 1'h0;
      end else begin
        mask_0_0_1 <= _GEN_1040;
      end
    end else begin
      mask_0_0_1 <= _GEN_1040;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_0_0_2 <= _GEN_8336;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_0_0_2 <= _GEN_4240; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_2 <= 1'h0;
      end else begin
        mask_0_0_2 <= _GEN_1056;
      end
    end else begin
      mask_0_0_2 <= _GEN_1056;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_0_0_3 <= _GEN_8400;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_0_0_3 <= _GEN_4304; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_3 <= 1'h0;
      end else begin
        mask_0_0_3 <= _GEN_1072;
      end
    end else begin
      mask_0_0_3 <= _GEN_1072;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_0_0_4 <= _GEN_8464;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_0_0_4 <= _GEN_4368; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_4 <= 1'h0;
      end else begin
        mask_0_0_4 <= _GEN_1088;
      end
    end else begin
      mask_0_0_4 <= _GEN_1088;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_0_0_5 <= _GEN_8528;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_0_0_5 <= _GEN_4432; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_5 <= 1'h0;
      end else begin
        mask_0_0_5 <= _GEN_1104;
      end
    end else begin
      mask_0_0_5 <= _GEN_1104;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_0_0_6 <= _GEN_8592;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_0_0_6 <= _GEN_4496; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_6 <= 1'h0;
      end else begin
        mask_0_0_6 <= _GEN_1120;
      end
    end else begin
      mask_0_0_6 <= _GEN_1120;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_0_0_7 <= _GEN_8656;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_0_0_7 <= _GEN_4560; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_0_7 <= 1'h0;
      end else begin
        mask_0_0_7 <= _GEN_1136;
      end
    end else begin
      mask_0_0_7 <= _GEN_1136;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_0_1_0 <= _GEN_8720;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_0_1_0 <= _GEN_4624; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_0 <= 1'h0;
      end else begin
        mask_0_1_0 <= _GEN_1152;
      end
    end else begin
      mask_0_1_0 <= _GEN_1152;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_0_1_1 <= _GEN_8784;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_0_1_1 <= _GEN_4688; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_1 <= 1'h0;
      end else begin
        mask_0_1_1 <= _GEN_1168;
      end
    end else begin
      mask_0_1_1 <= _GEN_1168;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_0_1_2 <= _GEN_8848;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_0_1_2 <= _GEN_4752; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_2 <= 1'h0;
      end else begin
        mask_0_1_2 <= _GEN_1184;
      end
    end else begin
      mask_0_1_2 <= _GEN_1184;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_0_1_3 <= _GEN_8912;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_0_1_3 <= _GEN_4816; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_3 <= 1'h0;
      end else begin
        mask_0_1_3 <= _GEN_1200;
      end
    end else begin
      mask_0_1_3 <= _GEN_1200;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_0_1_4 <= _GEN_8976;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_0_1_4 <= _GEN_4880; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_4 <= 1'h0;
      end else begin
        mask_0_1_4 <= _GEN_1216;
      end
    end else begin
      mask_0_1_4 <= _GEN_1216;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_0_1_5 <= _GEN_9040;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_0_1_5 <= _GEN_4944; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_5 <= 1'h0;
      end else begin
        mask_0_1_5 <= _GEN_1232;
      end
    end else begin
      mask_0_1_5 <= _GEN_1232;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_0_1_6 <= _GEN_9104;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_0_1_6 <= _GEN_5008; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_6 <= 1'h0;
      end else begin
        mask_0_1_6 <= _GEN_1248;
      end
    end else begin
      mask_0_1_6 <= _GEN_1248;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_0_1_7 <= _GEN_9168;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_0_1_7 <= _GEN_5072; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_1_7 <= 1'h0;
      end else begin
        mask_0_1_7 <= _GEN_1264;
      end
    end else begin
      mask_0_1_7 <= _GEN_1264;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_0_2_0 <= _GEN_9232;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_0_2_0 <= _GEN_5136; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_0 <= 1'h0;
      end else begin
        mask_0_2_0 <= _GEN_1280;
      end
    end else begin
      mask_0_2_0 <= _GEN_1280;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_0_2_1 <= _GEN_9296;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_0_2_1 <= _GEN_5200; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_1 <= 1'h0;
      end else begin
        mask_0_2_1 <= _GEN_1296;
      end
    end else begin
      mask_0_2_1 <= _GEN_1296;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_0_2_2 <= _GEN_9360;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_0_2_2 <= _GEN_5264; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_2 <= 1'h0;
      end else begin
        mask_0_2_2 <= _GEN_1312;
      end
    end else begin
      mask_0_2_2 <= _GEN_1312;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_0_2_3 <= _GEN_9424;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_0_2_3 <= _GEN_5328; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_3 <= 1'h0;
      end else begin
        mask_0_2_3 <= _GEN_1328;
      end
    end else begin
      mask_0_2_3 <= _GEN_1328;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_0_2_4 <= _GEN_9488;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_0_2_4 <= _GEN_5392; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_4 <= 1'h0;
      end else begin
        mask_0_2_4 <= _GEN_1344;
      end
    end else begin
      mask_0_2_4 <= _GEN_1344;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_0_2_5 <= _GEN_9552;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_0_2_5 <= _GEN_5456; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_5 <= 1'h0;
      end else begin
        mask_0_2_5 <= _GEN_1360;
      end
    end else begin
      mask_0_2_5 <= _GEN_1360;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_0_2_6 <= _GEN_9616;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_0_2_6 <= _GEN_5520; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_6 <= 1'h0;
      end else begin
        mask_0_2_6 <= _GEN_1376;
      end
    end else begin
      mask_0_2_6 <= _GEN_1376;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_0_2_7 <= _GEN_9680;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_0_2_7 <= _GEN_5584; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_2_7 <= 1'h0;
      end else begin
        mask_0_2_7 <= _GEN_1392;
      end
    end else begin
      mask_0_2_7 <= _GEN_1392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_0_3_0 <= _GEN_9744;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_0_3_0 <= _GEN_5648; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_0 <= 1'h0;
      end else begin
        mask_0_3_0 <= _GEN_1408;
      end
    end else begin
      mask_0_3_0 <= _GEN_1408;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_0_3_1 <= _GEN_9808;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_0_3_1 <= _GEN_5712; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_1 <= 1'h0;
      end else begin
        mask_0_3_1 <= _GEN_1424;
      end
    end else begin
      mask_0_3_1 <= _GEN_1424;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_0_3_2 <= _GEN_9872;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_0_3_2 <= _GEN_5776; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_2 <= 1'h0;
      end else begin
        mask_0_3_2 <= _GEN_1440;
      end
    end else begin
      mask_0_3_2 <= _GEN_1440;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_0_3_3 <= _GEN_9936;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_0_3_3 <= _GEN_5840; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_3 <= 1'h0;
      end else begin
        mask_0_3_3 <= _GEN_1456;
      end
    end else begin
      mask_0_3_3 <= _GEN_1456;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_0_3_4 <= _GEN_10000;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_0_3_4 <= _GEN_5904; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_4 <= 1'h0;
      end else begin
        mask_0_3_4 <= _GEN_1472;
      end
    end else begin
      mask_0_3_4 <= _GEN_1472;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_0_3_5 <= _GEN_10064;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_0_3_5 <= _GEN_5968; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_5 <= 1'h0;
      end else begin
        mask_0_3_5 <= _GEN_1488;
      end
    end else begin
      mask_0_3_5 <= _GEN_1488;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_0_3_6 <= _GEN_10128;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_0_3_6 <= _GEN_6032; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_6 <= 1'h0;
      end else begin
        mask_0_3_6 <= _GEN_1504;
      end
    end else begin
      mask_0_3_6 <= _GEN_1504;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_0_3_7 <= _GEN_10192;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_0_3_7 <= _GEN_6096; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_3_7 <= 1'h0;
      end else begin
        mask_0_3_7 <= _GEN_1520;
      end
    end else begin
      mask_0_3_7 <= _GEN_1520;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_0_4_0 <= _GEN_10256;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_0_4_0 <= _GEN_6160; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_0 <= 1'h0;
      end else begin
        mask_0_4_0 <= _GEN_1536;
      end
    end else begin
      mask_0_4_0 <= _GEN_1536;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_0_4_1 <= _GEN_10320;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_0_4_1 <= _GEN_6224; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_1 <= 1'h0;
      end else begin
        mask_0_4_1 <= _GEN_1552;
      end
    end else begin
      mask_0_4_1 <= _GEN_1552;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_0_4_2 <= _GEN_10384;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_0_4_2 <= _GEN_6288; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_2 <= 1'h0;
      end else begin
        mask_0_4_2 <= _GEN_1568;
      end
    end else begin
      mask_0_4_2 <= _GEN_1568;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_0_4_3 <= _GEN_10448;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_0_4_3 <= _GEN_6352; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_3 <= 1'h0;
      end else begin
        mask_0_4_3 <= _GEN_1584;
      end
    end else begin
      mask_0_4_3 <= _GEN_1584;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_0_4_4 <= _GEN_10512;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_0_4_4 <= _GEN_6416; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_4 <= 1'h0;
      end else begin
        mask_0_4_4 <= _GEN_1600;
      end
    end else begin
      mask_0_4_4 <= _GEN_1600;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_0_4_5 <= _GEN_10576;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_0_4_5 <= _GEN_6480; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_5 <= 1'h0;
      end else begin
        mask_0_4_5 <= _GEN_1616;
      end
    end else begin
      mask_0_4_5 <= _GEN_1616;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_0_4_6 <= _GEN_10640;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_0_4_6 <= _GEN_6544; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_6 <= 1'h0;
      end else begin
        mask_0_4_6 <= _GEN_1632;
      end
    end else begin
      mask_0_4_6 <= _GEN_1632;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_0_4_7 <= _GEN_10704;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_0_4_7 <= _GEN_6608; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_4_7 <= 1'h0;
      end else begin
        mask_0_4_7 <= _GEN_1648;
      end
    end else begin
      mask_0_4_7 <= _GEN_1648;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_0_5_0 <= _GEN_10768;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_0_5_0 <= _GEN_6672; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_0 <= 1'h0;
      end else begin
        mask_0_5_0 <= _GEN_1664;
      end
    end else begin
      mask_0_5_0 <= _GEN_1664;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_0_5_1 <= _GEN_10832;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_0_5_1 <= _GEN_6736; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_1 <= 1'h0;
      end else begin
        mask_0_5_1 <= _GEN_1680;
      end
    end else begin
      mask_0_5_1 <= _GEN_1680;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_0_5_2 <= _GEN_10896;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_0_5_2 <= _GEN_6800; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_2 <= 1'h0;
      end else begin
        mask_0_5_2 <= _GEN_1696;
      end
    end else begin
      mask_0_5_2 <= _GEN_1696;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_0_5_3 <= _GEN_10960;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_0_5_3 <= _GEN_6864; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_3 <= 1'h0;
      end else begin
        mask_0_5_3 <= _GEN_1712;
      end
    end else begin
      mask_0_5_3 <= _GEN_1712;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_0_5_4 <= _GEN_11024;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_0_5_4 <= _GEN_6928; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_4 <= 1'h0;
      end else begin
        mask_0_5_4 <= _GEN_1728;
      end
    end else begin
      mask_0_5_4 <= _GEN_1728;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_0_5_5 <= _GEN_11088;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_0_5_5 <= _GEN_6992; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_5 <= 1'h0;
      end else begin
        mask_0_5_5 <= _GEN_1744;
      end
    end else begin
      mask_0_5_5 <= _GEN_1744;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_0_5_6 <= _GEN_11152;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_0_5_6 <= _GEN_7056; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_6 <= 1'h0;
      end else begin
        mask_0_5_6 <= _GEN_1760;
      end
    end else begin
      mask_0_5_6 <= _GEN_1760;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_0_5_7 <= _GEN_11216;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_0_5_7 <= _GEN_7120; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_5_7 <= 1'h0;
      end else begin
        mask_0_5_7 <= _GEN_1776;
      end
    end else begin
      mask_0_5_7 <= _GEN_1776;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_0_6_0 <= _GEN_11280;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_0_6_0 <= _GEN_7184; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_0 <= 1'h0;
      end else begin
        mask_0_6_0 <= _GEN_1792;
      end
    end else begin
      mask_0_6_0 <= _GEN_1792;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_0_6_1 <= _GEN_11344;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_0_6_1 <= _GEN_7248; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_1 <= 1'h0;
      end else begin
        mask_0_6_1 <= _GEN_1808;
      end
    end else begin
      mask_0_6_1 <= _GEN_1808;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_0_6_2 <= _GEN_11408;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_0_6_2 <= _GEN_7312; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_2 <= 1'h0;
      end else begin
        mask_0_6_2 <= _GEN_1824;
      end
    end else begin
      mask_0_6_2 <= _GEN_1824;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_0_6_3 <= _GEN_11472;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_0_6_3 <= _GEN_7376; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_3 <= 1'h0;
      end else begin
        mask_0_6_3 <= _GEN_1840;
      end
    end else begin
      mask_0_6_3 <= _GEN_1840;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_0_6_4 <= _GEN_11536;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_0_6_4 <= _GEN_7440; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_4 <= 1'h0;
      end else begin
        mask_0_6_4 <= _GEN_1856;
      end
    end else begin
      mask_0_6_4 <= _GEN_1856;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_0_6_5 <= _GEN_11600;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_0_6_5 <= _GEN_7504; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_5 <= 1'h0;
      end else begin
        mask_0_6_5 <= _GEN_1872;
      end
    end else begin
      mask_0_6_5 <= _GEN_1872;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_0_6_6 <= _GEN_11664;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_0_6_6 <= _GEN_7568; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_6 <= 1'h0;
      end else begin
        mask_0_6_6 <= _GEN_1888;
      end
    end else begin
      mask_0_6_6 <= _GEN_1888;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_0_6_7 <= _GEN_11728;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_0_6_7 <= _GEN_7632; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_6_7 <= 1'h0;
      end else begin
        mask_0_6_7 <= _GEN_1904;
      end
    end else begin
      mask_0_6_7 <= _GEN_1904;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_0_7_0 <= _GEN_11792;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_0_7_0 <= _GEN_7696; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_0 <= 1'h0;
      end else begin
        mask_0_7_0 <= _GEN_1920;
      end
    end else begin
      mask_0_7_0 <= _GEN_1920;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_0_7_1 <= _GEN_11856;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_0_7_1 <= _GEN_7760; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_1 <= 1'h0;
      end else begin
        mask_0_7_1 <= _GEN_1936;
      end
    end else begin
      mask_0_7_1 <= _GEN_1936;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_0_7_2 <= _GEN_11920;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_0_7_2 <= _GEN_7824; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_2 <= 1'h0;
      end else begin
        mask_0_7_2 <= _GEN_1952;
      end
    end else begin
      mask_0_7_2 <= _GEN_1952;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_0_7_3 <= _GEN_11984;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_0_7_3 <= _GEN_7888; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_3 <= 1'h0;
      end else begin
        mask_0_7_3 <= _GEN_1968;
      end
    end else begin
      mask_0_7_3 <= _GEN_1968;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_0_7_4 <= _GEN_12048;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_0_7_4 <= _GEN_7952; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_4 <= 1'h0;
      end else begin
        mask_0_7_4 <= _GEN_1984;
      end
    end else begin
      mask_0_7_4 <= _GEN_1984;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_0_7_5 <= _GEN_12112;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_0_7_5 <= _GEN_8016; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_5 <= 1'h0;
      end else begin
        mask_0_7_5 <= _GEN_2000;
      end
    end else begin
      mask_0_7_5 <= _GEN_2000;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_0_7_6 <= _GEN_12176;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_0_7_6 <= _GEN_8080; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_6 <= 1'h0;
      end else begin
        mask_0_7_6 <= _GEN_2016;
      end
    end else begin
      mask_0_7_6 <= _GEN_2016;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_0_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_0_7_7 <= _GEN_12240;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_0_7_7 <= _GEN_8144; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h0 == line_mask_clean_line_1) begin
        mask_0_7_7 <= 1'h0;
      end else begin
        mask_0_7_7 <= _GEN_2032;
      end
    end else begin
      mask_0_7_7 <= _GEN_2032;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_1_0_0 <= _GEN_8209;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_1_0_0 <= _GEN_4113; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_0 <= 1'h0;
      end else begin
        mask_1_0_0 <= _GEN_1025;
      end
    end else begin
      mask_1_0_0 <= _GEN_1025;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_1_0_1 <= _GEN_8273;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_1_0_1 <= _GEN_4177; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_1 <= 1'h0;
      end else begin
        mask_1_0_1 <= _GEN_1041;
      end
    end else begin
      mask_1_0_1 <= _GEN_1041;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_1_0_2 <= _GEN_8337;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_1_0_2 <= _GEN_4241; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_2 <= 1'h0;
      end else begin
        mask_1_0_2 <= _GEN_1057;
      end
    end else begin
      mask_1_0_2 <= _GEN_1057;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_1_0_3 <= _GEN_8401;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_1_0_3 <= _GEN_4305; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_3 <= 1'h0;
      end else begin
        mask_1_0_3 <= _GEN_1073;
      end
    end else begin
      mask_1_0_3 <= _GEN_1073;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_1_0_4 <= _GEN_8465;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_1_0_4 <= _GEN_4369; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_4 <= 1'h0;
      end else begin
        mask_1_0_4 <= _GEN_1089;
      end
    end else begin
      mask_1_0_4 <= _GEN_1089;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_1_0_5 <= _GEN_8529;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_1_0_5 <= _GEN_4433; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_5 <= 1'h0;
      end else begin
        mask_1_0_5 <= _GEN_1105;
      end
    end else begin
      mask_1_0_5 <= _GEN_1105;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_1_0_6 <= _GEN_8593;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_1_0_6 <= _GEN_4497; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_6 <= 1'h0;
      end else begin
        mask_1_0_6 <= _GEN_1121;
      end
    end else begin
      mask_1_0_6 <= _GEN_1121;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_1_0_7 <= _GEN_8657;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_1_0_7 <= _GEN_4561; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_0_7 <= 1'h0;
      end else begin
        mask_1_0_7 <= _GEN_1137;
      end
    end else begin
      mask_1_0_7 <= _GEN_1137;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_1_1_0 <= _GEN_8721;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_1_1_0 <= _GEN_4625; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_0 <= 1'h0;
      end else begin
        mask_1_1_0 <= _GEN_1153;
      end
    end else begin
      mask_1_1_0 <= _GEN_1153;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_1_1_1 <= _GEN_8785;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_1_1_1 <= _GEN_4689; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_1 <= 1'h0;
      end else begin
        mask_1_1_1 <= _GEN_1169;
      end
    end else begin
      mask_1_1_1 <= _GEN_1169;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_1_1_2 <= _GEN_8849;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_1_1_2 <= _GEN_4753; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_2 <= 1'h0;
      end else begin
        mask_1_1_2 <= _GEN_1185;
      end
    end else begin
      mask_1_1_2 <= _GEN_1185;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_1_1_3 <= _GEN_8913;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_1_1_3 <= _GEN_4817; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_3 <= 1'h0;
      end else begin
        mask_1_1_3 <= _GEN_1201;
      end
    end else begin
      mask_1_1_3 <= _GEN_1201;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_1_1_4 <= _GEN_8977;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_1_1_4 <= _GEN_4881; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_4 <= 1'h0;
      end else begin
        mask_1_1_4 <= _GEN_1217;
      end
    end else begin
      mask_1_1_4 <= _GEN_1217;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_1_1_5 <= _GEN_9041;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_1_1_5 <= _GEN_4945; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_5 <= 1'h0;
      end else begin
        mask_1_1_5 <= _GEN_1233;
      end
    end else begin
      mask_1_1_5 <= _GEN_1233;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_1_1_6 <= _GEN_9105;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_1_1_6 <= _GEN_5009; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_6 <= 1'h0;
      end else begin
        mask_1_1_6 <= _GEN_1249;
      end
    end else begin
      mask_1_1_6 <= _GEN_1249;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_1_1_7 <= _GEN_9169;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_1_1_7 <= _GEN_5073; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_1_7 <= 1'h0;
      end else begin
        mask_1_1_7 <= _GEN_1265;
      end
    end else begin
      mask_1_1_7 <= _GEN_1265;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_1_2_0 <= _GEN_9233;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_1_2_0 <= _GEN_5137; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_0 <= 1'h0;
      end else begin
        mask_1_2_0 <= _GEN_1281;
      end
    end else begin
      mask_1_2_0 <= _GEN_1281;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_1_2_1 <= _GEN_9297;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_1_2_1 <= _GEN_5201; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_1 <= 1'h0;
      end else begin
        mask_1_2_1 <= _GEN_1297;
      end
    end else begin
      mask_1_2_1 <= _GEN_1297;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_1_2_2 <= _GEN_9361;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_1_2_2 <= _GEN_5265; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_2 <= 1'h0;
      end else begin
        mask_1_2_2 <= _GEN_1313;
      end
    end else begin
      mask_1_2_2 <= _GEN_1313;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_1_2_3 <= _GEN_9425;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_1_2_3 <= _GEN_5329; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_3 <= 1'h0;
      end else begin
        mask_1_2_3 <= _GEN_1329;
      end
    end else begin
      mask_1_2_3 <= _GEN_1329;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_1_2_4 <= _GEN_9489;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_1_2_4 <= _GEN_5393; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_4 <= 1'h0;
      end else begin
        mask_1_2_4 <= _GEN_1345;
      end
    end else begin
      mask_1_2_4 <= _GEN_1345;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_1_2_5 <= _GEN_9553;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_1_2_5 <= _GEN_5457; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_5 <= 1'h0;
      end else begin
        mask_1_2_5 <= _GEN_1361;
      end
    end else begin
      mask_1_2_5 <= _GEN_1361;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_1_2_6 <= _GEN_9617;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_1_2_6 <= _GEN_5521; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_6 <= 1'h0;
      end else begin
        mask_1_2_6 <= _GEN_1377;
      end
    end else begin
      mask_1_2_6 <= _GEN_1377;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_1_2_7 <= _GEN_9681;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_1_2_7 <= _GEN_5585; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_2_7 <= 1'h0;
      end else begin
        mask_1_2_7 <= _GEN_1393;
      end
    end else begin
      mask_1_2_7 <= _GEN_1393;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_1_3_0 <= _GEN_9745;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_1_3_0 <= _GEN_5649; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_0 <= 1'h0;
      end else begin
        mask_1_3_0 <= _GEN_1409;
      end
    end else begin
      mask_1_3_0 <= _GEN_1409;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_1_3_1 <= _GEN_9809;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_1_3_1 <= _GEN_5713; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_1 <= 1'h0;
      end else begin
        mask_1_3_1 <= _GEN_1425;
      end
    end else begin
      mask_1_3_1 <= _GEN_1425;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_1_3_2 <= _GEN_9873;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_1_3_2 <= _GEN_5777; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_2 <= 1'h0;
      end else begin
        mask_1_3_2 <= _GEN_1441;
      end
    end else begin
      mask_1_3_2 <= _GEN_1441;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_1_3_3 <= _GEN_9937;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_1_3_3 <= _GEN_5841; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_3 <= 1'h0;
      end else begin
        mask_1_3_3 <= _GEN_1457;
      end
    end else begin
      mask_1_3_3 <= _GEN_1457;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_1_3_4 <= _GEN_10001;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_1_3_4 <= _GEN_5905; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_4 <= 1'h0;
      end else begin
        mask_1_3_4 <= _GEN_1473;
      end
    end else begin
      mask_1_3_4 <= _GEN_1473;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_1_3_5 <= _GEN_10065;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_1_3_5 <= _GEN_5969; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_5 <= 1'h0;
      end else begin
        mask_1_3_5 <= _GEN_1489;
      end
    end else begin
      mask_1_3_5 <= _GEN_1489;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_1_3_6 <= _GEN_10129;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_1_3_6 <= _GEN_6033; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_6 <= 1'h0;
      end else begin
        mask_1_3_6 <= _GEN_1505;
      end
    end else begin
      mask_1_3_6 <= _GEN_1505;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_1_3_7 <= _GEN_10193;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_1_3_7 <= _GEN_6097; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_3_7 <= 1'h0;
      end else begin
        mask_1_3_7 <= _GEN_1521;
      end
    end else begin
      mask_1_3_7 <= _GEN_1521;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_1_4_0 <= _GEN_10257;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_1_4_0 <= _GEN_6161; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_0 <= 1'h0;
      end else begin
        mask_1_4_0 <= _GEN_1537;
      end
    end else begin
      mask_1_4_0 <= _GEN_1537;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_1_4_1 <= _GEN_10321;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_1_4_1 <= _GEN_6225; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_1 <= 1'h0;
      end else begin
        mask_1_4_1 <= _GEN_1553;
      end
    end else begin
      mask_1_4_1 <= _GEN_1553;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_1_4_2 <= _GEN_10385;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_1_4_2 <= _GEN_6289; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_2 <= 1'h0;
      end else begin
        mask_1_4_2 <= _GEN_1569;
      end
    end else begin
      mask_1_4_2 <= _GEN_1569;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_1_4_3 <= _GEN_10449;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_1_4_3 <= _GEN_6353; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_3 <= 1'h0;
      end else begin
        mask_1_4_3 <= _GEN_1585;
      end
    end else begin
      mask_1_4_3 <= _GEN_1585;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_1_4_4 <= _GEN_10513;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_1_4_4 <= _GEN_6417; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_4 <= 1'h0;
      end else begin
        mask_1_4_4 <= _GEN_1601;
      end
    end else begin
      mask_1_4_4 <= _GEN_1601;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_1_4_5 <= _GEN_10577;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_1_4_5 <= _GEN_6481; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_5 <= 1'h0;
      end else begin
        mask_1_4_5 <= _GEN_1617;
      end
    end else begin
      mask_1_4_5 <= _GEN_1617;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_1_4_6 <= _GEN_10641;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_1_4_6 <= _GEN_6545; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_6 <= 1'h0;
      end else begin
        mask_1_4_6 <= _GEN_1633;
      end
    end else begin
      mask_1_4_6 <= _GEN_1633;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_1_4_7 <= _GEN_10705;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_1_4_7 <= _GEN_6609; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_4_7 <= 1'h0;
      end else begin
        mask_1_4_7 <= _GEN_1649;
      end
    end else begin
      mask_1_4_7 <= _GEN_1649;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_1_5_0 <= _GEN_10769;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_1_5_0 <= _GEN_6673; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_0 <= 1'h0;
      end else begin
        mask_1_5_0 <= _GEN_1665;
      end
    end else begin
      mask_1_5_0 <= _GEN_1665;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_1_5_1 <= _GEN_10833;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_1_5_1 <= _GEN_6737; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_1 <= 1'h0;
      end else begin
        mask_1_5_1 <= _GEN_1681;
      end
    end else begin
      mask_1_5_1 <= _GEN_1681;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_1_5_2 <= _GEN_10897;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_1_5_2 <= _GEN_6801; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_2 <= 1'h0;
      end else begin
        mask_1_5_2 <= _GEN_1697;
      end
    end else begin
      mask_1_5_2 <= _GEN_1697;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_1_5_3 <= _GEN_10961;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_1_5_3 <= _GEN_6865; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_3 <= 1'h0;
      end else begin
        mask_1_5_3 <= _GEN_1713;
      end
    end else begin
      mask_1_5_3 <= _GEN_1713;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_1_5_4 <= _GEN_11025;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_1_5_4 <= _GEN_6929; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_4 <= 1'h0;
      end else begin
        mask_1_5_4 <= _GEN_1729;
      end
    end else begin
      mask_1_5_4 <= _GEN_1729;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_1_5_5 <= _GEN_11089;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_1_5_5 <= _GEN_6993; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_5 <= 1'h0;
      end else begin
        mask_1_5_5 <= _GEN_1745;
      end
    end else begin
      mask_1_5_5 <= _GEN_1745;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_1_5_6 <= _GEN_11153;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_1_5_6 <= _GEN_7057; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_6 <= 1'h0;
      end else begin
        mask_1_5_6 <= _GEN_1761;
      end
    end else begin
      mask_1_5_6 <= _GEN_1761;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_1_5_7 <= _GEN_11217;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_1_5_7 <= _GEN_7121; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_5_7 <= 1'h0;
      end else begin
        mask_1_5_7 <= _GEN_1777;
      end
    end else begin
      mask_1_5_7 <= _GEN_1777;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_1_6_0 <= _GEN_11281;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_1_6_0 <= _GEN_7185; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_0 <= 1'h0;
      end else begin
        mask_1_6_0 <= _GEN_1793;
      end
    end else begin
      mask_1_6_0 <= _GEN_1793;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_1_6_1 <= _GEN_11345;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_1_6_1 <= _GEN_7249; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_1 <= 1'h0;
      end else begin
        mask_1_6_1 <= _GEN_1809;
      end
    end else begin
      mask_1_6_1 <= _GEN_1809;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_1_6_2 <= _GEN_11409;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_1_6_2 <= _GEN_7313; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_2 <= 1'h0;
      end else begin
        mask_1_6_2 <= _GEN_1825;
      end
    end else begin
      mask_1_6_2 <= _GEN_1825;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_1_6_3 <= _GEN_11473;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_1_6_3 <= _GEN_7377; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_3 <= 1'h0;
      end else begin
        mask_1_6_3 <= _GEN_1841;
      end
    end else begin
      mask_1_6_3 <= _GEN_1841;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_1_6_4 <= _GEN_11537;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_1_6_4 <= _GEN_7441; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_4 <= 1'h0;
      end else begin
        mask_1_6_4 <= _GEN_1857;
      end
    end else begin
      mask_1_6_4 <= _GEN_1857;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_1_6_5 <= _GEN_11601;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_1_6_5 <= _GEN_7505; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_5 <= 1'h0;
      end else begin
        mask_1_6_5 <= _GEN_1873;
      end
    end else begin
      mask_1_6_5 <= _GEN_1873;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_1_6_6 <= _GEN_11665;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_1_6_6 <= _GEN_7569; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_6 <= 1'h0;
      end else begin
        mask_1_6_6 <= _GEN_1889;
      end
    end else begin
      mask_1_6_6 <= _GEN_1889;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_1_6_7 <= _GEN_11729;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_1_6_7 <= _GEN_7633; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_6_7 <= 1'h0;
      end else begin
        mask_1_6_7 <= _GEN_1905;
      end
    end else begin
      mask_1_6_7 <= _GEN_1905;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_1_7_0 <= _GEN_11793;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_1_7_0 <= _GEN_7697; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_0 <= 1'h0;
      end else begin
        mask_1_7_0 <= _GEN_1921;
      end
    end else begin
      mask_1_7_0 <= _GEN_1921;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_1_7_1 <= _GEN_11857;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_1_7_1 <= _GEN_7761; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_1 <= 1'h0;
      end else begin
        mask_1_7_1 <= _GEN_1937;
      end
    end else begin
      mask_1_7_1 <= _GEN_1937;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_1_7_2 <= _GEN_11921;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_1_7_2 <= _GEN_7825; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_2 <= 1'h0;
      end else begin
        mask_1_7_2 <= _GEN_1953;
      end
    end else begin
      mask_1_7_2 <= _GEN_1953;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_1_7_3 <= _GEN_11985;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_1_7_3 <= _GEN_7889; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_3 <= 1'h0;
      end else begin
        mask_1_7_3 <= _GEN_1969;
      end
    end else begin
      mask_1_7_3 <= _GEN_1969;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_1_7_4 <= _GEN_12049;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_1_7_4 <= _GEN_7953; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_4 <= 1'h0;
      end else begin
        mask_1_7_4 <= _GEN_1985;
      end
    end else begin
      mask_1_7_4 <= _GEN_1985;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_1_7_5 <= _GEN_12113;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_1_7_5 <= _GEN_8017; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_5 <= 1'h0;
      end else begin
        mask_1_7_5 <= _GEN_2001;
      end
    end else begin
      mask_1_7_5 <= _GEN_2001;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_1_7_6 <= _GEN_12177;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_1_7_6 <= _GEN_8081; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_6 <= 1'h0;
      end else begin
        mask_1_7_6 <= _GEN_2017;
      end
    end else begin
      mask_1_7_6 <= _GEN_2017;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_1_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_1_7_7 <= _GEN_12241;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_1_7_7 <= _GEN_8145; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h1 == line_mask_clean_line_1) begin
        mask_1_7_7 <= 1'h0;
      end else begin
        mask_1_7_7 <= _GEN_2033;
      end
    end else begin
      mask_1_7_7 <= _GEN_2033;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_2_0_0 <= _GEN_8210;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_2_0_0 <= _GEN_4114; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_0 <= 1'h0;
      end else begin
        mask_2_0_0 <= _GEN_1026;
      end
    end else begin
      mask_2_0_0 <= _GEN_1026;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_2_0_1 <= _GEN_8274;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_2_0_1 <= _GEN_4178; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_1 <= 1'h0;
      end else begin
        mask_2_0_1 <= _GEN_1042;
      end
    end else begin
      mask_2_0_1 <= _GEN_1042;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_2_0_2 <= _GEN_8338;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_2_0_2 <= _GEN_4242; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_2 <= 1'h0;
      end else begin
        mask_2_0_2 <= _GEN_1058;
      end
    end else begin
      mask_2_0_2 <= _GEN_1058;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_2_0_3 <= _GEN_8402;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_2_0_3 <= _GEN_4306; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_3 <= 1'h0;
      end else begin
        mask_2_0_3 <= _GEN_1074;
      end
    end else begin
      mask_2_0_3 <= _GEN_1074;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_2_0_4 <= _GEN_8466;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_2_0_4 <= _GEN_4370; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_4 <= 1'h0;
      end else begin
        mask_2_0_4 <= _GEN_1090;
      end
    end else begin
      mask_2_0_4 <= _GEN_1090;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_2_0_5 <= _GEN_8530;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_2_0_5 <= _GEN_4434; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_5 <= 1'h0;
      end else begin
        mask_2_0_5 <= _GEN_1106;
      end
    end else begin
      mask_2_0_5 <= _GEN_1106;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_2_0_6 <= _GEN_8594;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_2_0_6 <= _GEN_4498; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_6 <= 1'h0;
      end else begin
        mask_2_0_6 <= _GEN_1122;
      end
    end else begin
      mask_2_0_6 <= _GEN_1122;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_2_0_7 <= _GEN_8658;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_2_0_7 <= _GEN_4562; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_0_7 <= 1'h0;
      end else begin
        mask_2_0_7 <= _GEN_1138;
      end
    end else begin
      mask_2_0_7 <= _GEN_1138;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_2_1_0 <= _GEN_8722;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_2_1_0 <= _GEN_4626; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_0 <= 1'h0;
      end else begin
        mask_2_1_0 <= _GEN_1154;
      end
    end else begin
      mask_2_1_0 <= _GEN_1154;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_2_1_1 <= _GEN_8786;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_2_1_1 <= _GEN_4690; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_1 <= 1'h0;
      end else begin
        mask_2_1_1 <= _GEN_1170;
      end
    end else begin
      mask_2_1_1 <= _GEN_1170;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_2_1_2 <= _GEN_8850;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_2_1_2 <= _GEN_4754; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_2 <= 1'h0;
      end else begin
        mask_2_1_2 <= _GEN_1186;
      end
    end else begin
      mask_2_1_2 <= _GEN_1186;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_2_1_3 <= _GEN_8914;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_2_1_3 <= _GEN_4818; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_3 <= 1'h0;
      end else begin
        mask_2_1_3 <= _GEN_1202;
      end
    end else begin
      mask_2_1_3 <= _GEN_1202;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_2_1_4 <= _GEN_8978;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_2_1_4 <= _GEN_4882; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_4 <= 1'h0;
      end else begin
        mask_2_1_4 <= _GEN_1218;
      end
    end else begin
      mask_2_1_4 <= _GEN_1218;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_2_1_5 <= _GEN_9042;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_2_1_5 <= _GEN_4946; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_5 <= 1'h0;
      end else begin
        mask_2_1_5 <= _GEN_1234;
      end
    end else begin
      mask_2_1_5 <= _GEN_1234;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_2_1_6 <= _GEN_9106;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_2_1_6 <= _GEN_5010; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_6 <= 1'h0;
      end else begin
        mask_2_1_6 <= _GEN_1250;
      end
    end else begin
      mask_2_1_6 <= _GEN_1250;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_2_1_7 <= _GEN_9170;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_2_1_7 <= _GEN_5074; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_1_7 <= 1'h0;
      end else begin
        mask_2_1_7 <= _GEN_1266;
      end
    end else begin
      mask_2_1_7 <= _GEN_1266;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_2_2_0 <= _GEN_9234;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_2_2_0 <= _GEN_5138; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_0 <= 1'h0;
      end else begin
        mask_2_2_0 <= _GEN_1282;
      end
    end else begin
      mask_2_2_0 <= _GEN_1282;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_2_2_1 <= _GEN_9298;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_2_2_1 <= _GEN_5202; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_1 <= 1'h0;
      end else begin
        mask_2_2_1 <= _GEN_1298;
      end
    end else begin
      mask_2_2_1 <= _GEN_1298;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_2_2_2 <= _GEN_9362;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_2_2_2 <= _GEN_5266; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_2 <= 1'h0;
      end else begin
        mask_2_2_2 <= _GEN_1314;
      end
    end else begin
      mask_2_2_2 <= _GEN_1314;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_2_2_3 <= _GEN_9426;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_2_2_3 <= _GEN_5330; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_3 <= 1'h0;
      end else begin
        mask_2_2_3 <= _GEN_1330;
      end
    end else begin
      mask_2_2_3 <= _GEN_1330;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_2_2_4 <= _GEN_9490;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_2_2_4 <= _GEN_5394; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_4 <= 1'h0;
      end else begin
        mask_2_2_4 <= _GEN_1346;
      end
    end else begin
      mask_2_2_4 <= _GEN_1346;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_2_2_5 <= _GEN_9554;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_2_2_5 <= _GEN_5458; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_5 <= 1'h0;
      end else begin
        mask_2_2_5 <= _GEN_1362;
      end
    end else begin
      mask_2_2_5 <= _GEN_1362;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_2_2_6 <= _GEN_9618;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_2_2_6 <= _GEN_5522; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_6 <= 1'h0;
      end else begin
        mask_2_2_6 <= _GEN_1378;
      end
    end else begin
      mask_2_2_6 <= _GEN_1378;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_2_2_7 <= _GEN_9682;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_2_2_7 <= _GEN_5586; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_2_7 <= 1'h0;
      end else begin
        mask_2_2_7 <= _GEN_1394;
      end
    end else begin
      mask_2_2_7 <= _GEN_1394;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_2_3_0 <= _GEN_9746;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_2_3_0 <= _GEN_5650; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_0 <= 1'h0;
      end else begin
        mask_2_3_0 <= _GEN_1410;
      end
    end else begin
      mask_2_3_0 <= _GEN_1410;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_2_3_1 <= _GEN_9810;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_2_3_1 <= _GEN_5714; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_1 <= 1'h0;
      end else begin
        mask_2_3_1 <= _GEN_1426;
      end
    end else begin
      mask_2_3_1 <= _GEN_1426;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_2_3_2 <= _GEN_9874;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_2_3_2 <= _GEN_5778; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_2 <= 1'h0;
      end else begin
        mask_2_3_2 <= _GEN_1442;
      end
    end else begin
      mask_2_3_2 <= _GEN_1442;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_2_3_3 <= _GEN_9938;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_2_3_3 <= _GEN_5842; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_3 <= 1'h0;
      end else begin
        mask_2_3_3 <= _GEN_1458;
      end
    end else begin
      mask_2_3_3 <= _GEN_1458;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_2_3_4 <= _GEN_10002;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_2_3_4 <= _GEN_5906; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_4 <= 1'h0;
      end else begin
        mask_2_3_4 <= _GEN_1474;
      end
    end else begin
      mask_2_3_4 <= _GEN_1474;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_2_3_5 <= _GEN_10066;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_2_3_5 <= _GEN_5970; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_5 <= 1'h0;
      end else begin
        mask_2_3_5 <= _GEN_1490;
      end
    end else begin
      mask_2_3_5 <= _GEN_1490;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_2_3_6 <= _GEN_10130;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_2_3_6 <= _GEN_6034; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_6 <= 1'h0;
      end else begin
        mask_2_3_6 <= _GEN_1506;
      end
    end else begin
      mask_2_3_6 <= _GEN_1506;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_2_3_7 <= _GEN_10194;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_2_3_7 <= _GEN_6098; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_3_7 <= 1'h0;
      end else begin
        mask_2_3_7 <= _GEN_1522;
      end
    end else begin
      mask_2_3_7 <= _GEN_1522;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_2_4_0 <= _GEN_10258;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_2_4_0 <= _GEN_6162; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_0 <= 1'h0;
      end else begin
        mask_2_4_0 <= _GEN_1538;
      end
    end else begin
      mask_2_4_0 <= _GEN_1538;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_2_4_1 <= _GEN_10322;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_2_4_1 <= _GEN_6226; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_1 <= 1'h0;
      end else begin
        mask_2_4_1 <= _GEN_1554;
      end
    end else begin
      mask_2_4_1 <= _GEN_1554;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_2_4_2 <= _GEN_10386;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_2_4_2 <= _GEN_6290; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_2 <= 1'h0;
      end else begin
        mask_2_4_2 <= _GEN_1570;
      end
    end else begin
      mask_2_4_2 <= _GEN_1570;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_2_4_3 <= _GEN_10450;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_2_4_3 <= _GEN_6354; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_3 <= 1'h0;
      end else begin
        mask_2_4_3 <= _GEN_1586;
      end
    end else begin
      mask_2_4_3 <= _GEN_1586;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_2_4_4 <= _GEN_10514;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_2_4_4 <= _GEN_6418; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_4 <= 1'h0;
      end else begin
        mask_2_4_4 <= _GEN_1602;
      end
    end else begin
      mask_2_4_4 <= _GEN_1602;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_2_4_5 <= _GEN_10578;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_2_4_5 <= _GEN_6482; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_5 <= 1'h0;
      end else begin
        mask_2_4_5 <= _GEN_1618;
      end
    end else begin
      mask_2_4_5 <= _GEN_1618;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_2_4_6 <= _GEN_10642;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_2_4_6 <= _GEN_6546; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_6 <= 1'h0;
      end else begin
        mask_2_4_6 <= _GEN_1634;
      end
    end else begin
      mask_2_4_6 <= _GEN_1634;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_2_4_7 <= _GEN_10706;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_2_4_7 <= _GEN_6610; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_4_7 <= 1'h0;
      end else begin
        mask_2_4_7 <= _GEN_1650;
      end
    end else begin
      mask_2_4_7 <= _GEN_1650;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_2_5_0 <= _GEN_10770;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_2_5_0 <= _GEN_6674; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_0 <= 1'h0;
      end else begin
        mask_2_5_0 <= _GEN_1666;
      end
    end else begin
      mask_2_5_0 <= _GEN_1666;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_2_5_1 <= _GEN_10834;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_2_5_1 <= _GEN_6738; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_1 <= 1'h0;
      end else begin
        mask_2_5_1 <= _GEN_1682;
      end
    end else begin
      mask_2_5_1 <= _GEN_1682;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_2_5_2 <= _GEN_10898;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_2_5_2 <= _GEN_6802; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_2 <= 1'h0;
      end else begin
        mask_2_5_2 <= _GEN_1698;
      end
    end else begin
      mask_2_5_2 <= _GEN_1698;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_2_5_3 <= _GEN_10962;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_2_5_3 <= _GEN_6866; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_3 <= 1'h0;
      end else begin
        mask_2_5_3 <= _GEN_1714;
      end
    end else begin
      mask_2_5_3 <= _GEN_1714;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_2_5_4 <= _GEN_11026;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_2_5_4 <= _GEN_6930; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_4 <= 1'h0;
      end else begin
        mask_2_5_4 <= _GEN_1730;
      end
    end else begin
      mask_2_5_4 <= _GEN_1730;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_2_5_5 <= _GEN_11090;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_2_5_5 <= _GEN_6994; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_5 <= 1'h0;
      end else begin
        mask_2_5_5 <= _GEN_1746;
      end
    end else begin
      mask_2_5_5 <= _GEN_1746;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_2_5_6 <= _GEN_11154;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_2_5_6 <= _GEN_7058; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_6 <= 1'h0;
      end else begin
        mask_2_5_6 <= _GEN_1762;
      end
    end else begin
      mask_2_5_6 <= _GEN_1762;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_2_5_7 <= _GEN_11218;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_2_5_7 <= _GEN_7122; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_5_7 <= 1'h0;
      end else begin
        mask_2_5_7 <= _GEN_1778;
      end
    end else begin
      mask_2_5_7 <= _GEN_1778;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_2_6_0 <= _GEN_11282;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_2_6_0 <= _GEN_7186; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_0 <= 1'h0;
      end else begin
        mask_2_6_0 <= _GEN_1794;
      end
    end else begin
      mask_2_6_0 <= _GEN_1794;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_2_6_1 <= _GEN_11346;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_2_6_1 <= _GEN_7250; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_1 <= 1'h0;
      end else begin
        mask_2_6_1 <= _GEN_1810;
      end
    end else begin
      mask_2_6_1 <= _GEN_1810;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_2_6_2 <= _GEN_11410;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_2_6_2 <= _GEN_7314; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_2 <= 1'h0;
      end else begin
        mask_2_6_2 <= _GEN_1826;
      end
    end else begin
      mask_2_6_2 <= _GEN_1826;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_2_6_3 <= _GEN_11474;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_2_6_3 <= _GEN_7378; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_3 <= 1'h0;
      end else begin
        mask_2_6_3 <= _GEN_1842;
      end
    end else begin
      mask_2_6_3 <= _GEN_1842;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_2_6_4 <= _GEN_11538;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_2_6_4 <= _GEN_7442; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_4 <= 1'h0;
      end else begin
        mask_2_6_4 <= _GEN_1858;
      end
    end else begin
      mask_2_6_4 <= _GEN_1858;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_2_6_5 <= _GEN_11602;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_2_6_5 <= _GEN_7506; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_5 <= 1'h0;
      end else begin
        mask_2_6_5 <= _GEN_1874;
      end
    end else begin
      mask_2_6_5 <= _GEN_1874;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_2_6_6 <= _GEN_11666;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_2_6_6 <= _GEN_7570; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_6 <= 1'h0;
      end else begin
        mask_2_6_6 <= _GEN_1890;
      end
    end else begin
      mask_2_6_6 <= _GEN_1890;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_2_6_7 <= _GEN_11730;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_2_6_7 <= _GEN_7634; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_6_7 <= 1'h0;
      end else begin
        mask_2_6_7 <= _GEN_1906;
      end
    end else begin
      mask_2_6_7 <= _GEN_1906;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_2_7_0 <= _GEN_11794;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_2_7_0 <= _GEN_7698; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_0 <= 1'h0;
      end else begin
        mask_2_7_0 <= _GEN_1922;
      end
    end else begin
      mask_2_7_0 <= _GEN_1922;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_2_7_1 <= _GEN_11858;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_2_7_1 <= _GEN_7762; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_1 <= 1'h0;
      end else begin
        mask_2_7_1 <= _GEN_1938;
      end
    end else begin
      mask_2_7_1 <= _GEN_1938;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_2_7_2 <= _GEN_11922;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_2_7_2 <= _GEN_7826; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_2 <= 1'h0;
      end else begin
        mask_2_7_2 <= _GEN_1954;
      end
    end else begin
      mask_2_7_2 <= _GEN_1954;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_2_7_3 <= _GEN_11986;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_2_7_3 <= _GEN_7890; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_3 <= 1'h0;
      end else begin
        mask_2_7_3 <= _GEN_1970;
      end
    end else begin
      mask_2_7_3 <= _GEN_1970;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_2_7_4 <= _GEN_12050;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_2_7_4 <= _GEN_7954; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_4 <= 1'h0;
      end else begin
        mask_2_7_4 <= _GEN_1986;
      end
    end else begin
      mask_2_7_4 <= _GEN_1986;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_2_7_5 <= _GEN_12114;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_2_7_5 <= _GEN_8018; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_5 <= 1'h0;
      end else begin
        mask_2_7_5 <= _GEN_2002;
      end
    end else begin
      mask_2_7_5 <= _GEN_2002;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_2_7_6 <= _GEN_12178;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_2_7_6 <= _GEN_8082; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_6 <= 1'h0;
      end else begin
        mask_2_7_6 <= _GEN_2018;
      end
    end else begin
      mask_2_7_6 <= _GEN_2018;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_2_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_2_7_7 <= _GEN_12242;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_2_7_7 <= _GEN_8146; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h2 == line_mask_clean_line_1) begin
        mask_2_7_7 <= 1'h0;
      end else begin
        mask_2_7_7 <= _GEN_2034;
      end
    end else begin
      mask_2_7_7 <= _GEN_2034;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_3_0_0 <= _GEN_8211;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_3_0_0 <= _GEN_4115; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_0 <= 1'h0;
      end else begin
        mask_3_0_0 <= _GEN_1027;
      end
    end else begin
      mask_3_0_0 <= _GEN_1027;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_3_0_1 <= _GEN_8275;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_3_0_1 <= _GEN_4179; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_1 <= 1'h0;
      end else begin
        mask_3_0_1 <= _GEN_1043;
      end
    end else begin
      mask_3_0_1 <= _GEN_1043;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_3_0_2 <= _GEN_8339;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_3_0_2 <= _GEN_4243; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_2 <= 1'h0;
      end else begin
        mask_3_0_2 <= _GEN_1059;
      end
    end else begin
      mask_3_0_2 <= _GEN_1059;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_3_0_3 <= _GEN_8403;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_3_0_3 <= _GEN_4307; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_3 <= 1'h0;
      end else begin
        mask_3_0_3 <= _GEN_1075;
      end
    end else begin
      mask_3_0_3 <= _GEN_1075;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_3_0_4 <= _GEN_8467;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_3_0_4 <= _GEN_4371; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_4 <= 1'h0;
      end else begin
        mask_3_0_4 <= _GEN_1091;
      end
    end else begin
      mask_3_0_4 <= _GEN_1091;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_3_0_5 <= _GEN_8531;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_3_0_5 <= _GEN_4435; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_5 <= 1'h0;
      end else begin
        mask_3_0_5 <= _GEN_1107;
      end
    end else begin
      mask_3_0_5 <= _GEN_1107;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_3_0_6 <= _GEN_8595;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_3_0_6 <= _GEN_4499; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_6 <= 1'h0;
      end else begin
        mask_3_0_6 <= _GEN_1123;
      end
    end else begin
      mask_3_0_6 <= _GEN_1123;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_3_0_7 <= _GEN_8659;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_3_0_7 <= _GEN_4563; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_0_7 <= 1'h0;
      end else begin
        mask_3_0_7 <= _GEN_1139;
      end
    end else begin
      mask_3_0_7 <= _GEN_1139;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_3_1_0 <= _GEN_8723;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_3_1_0 <= _GEN_4627; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_0 <= 1'h0;
      end else begin
        mask_3_1_0 <= _GEN_1155;
      end
    end else begin
      mask_3_1_0 <= _GEN_1155;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_3_1_1 <= _GEN_8787;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_3_1_1 <= _GEN_4691; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_1 <= 1'h0;
      end else begin
        mask_3_1_1 <= _GEN_1171;
      end
    end else begin
      mask_3_1_1 <= _GEN_1171;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_3_1_2 <= _GEN_8851;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_3_1_2 <= _GEN_4755; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_2 <= 1'h0;
      end else begin
        mask_3_1_2 <= _GEN_1187;
      end
    end else begin
      mask_3_1_2 <= _GEN_1187;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_3_1_3 <= _GEN_8915;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_3_1_3 <= _GEN_4819; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_3 <= 1'h0;
      end else begin
        mask_3_1_3 <= _GEN_1203;
      end
    end else begin
      mask_3_1_3 <= _GEN_1203;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_3_1_4 <= _GEN_8979;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_3_1_4 <= _GEN_4883; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_4 <= 1'h0;
      end else begin
        mask_3_1_4 <= _GEN_1219;
      end
    end else begin
      mask_3_1_4 <= _GEN_1219;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_3_1_5 <= _GEN_9043;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_3_1_5 <= _GEN_4947; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_5 <= 1'h0;
      end else begin
        mask_3_1_5 <= _GEN_1235;
      end
    end else begin
      mask_3_1_5 <= _GEN_1235;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_3_1_6 <= _GEN_9107;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_3_1_6 <= _GEN_5011; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_6 <= 1'h0;
      end else begin
        mask_3_1_6 <= _GEN_1251;
      end
    end else begin
      mask_3_1_6 <= _GEN_1251;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_3_1_7 <= _GEN_9171;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_3_1_7 <= _GEN_5075; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_1_7 <= 1'h0;
      end else begin
        mask_3_1_7 <= _GEN_1267;
      end
    end else begin
      mask_3_1_7 <= _GEN_1267;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_3_2_0 <= _GEN_9235;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_3_2_0 <= _GEN_5139; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_0 <= 1'h0;
      end else begin
        mask_3_2_0 <= _GEN_1283;
      end
    end else begin
      mask_3_2_0 <= _GEN_1283;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_3_2_1 <= _GEN_9299;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_3_2_1 <= _GEN_5203; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_1 <= 1'h0;
      end else begin
        mask_3_2_1 <= _GEN_1299;
      end
    end else begin
      mask_3_2_1 <= _GEN_1299;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_3_2_2 <= _GEN_9363;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_3_2_2 <= _GEN_5267; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_2 <= 1'h0;
      end else begin
        mask_3_2_2 <= _GEN_1315;
      end
    end else begin
      mask_3_2_2 <= _GEN_1315;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_3_2_3 <= _GEN_9427;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_3_2_3 <= _GEN_5331; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_3 <= 1'h0;
      end else begin
        mask_3_2_3 <= _GEN_1331;
      end
    end else begin
      mask_3_2_3 <= _GEN_1331;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_3_2_4 <= _GEN_9491;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_3_2_4 <= _GEN_5395; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_4 <= 1'h0;
      end else begin
        mask_3_2_4 <= _GEN_1347;
      end
    end else begin
      mask_3_2_4 <= _GEN_1347;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_3_2_5 <= _GEN_9555;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_3_2_5 <= _GEN_5459; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_5 <= 1'h0;
      end else begin
        mask_3_2_5 <= _GEN_1363;
      end
    end else begin
      mask_3_2_5 <= _GEN_1363;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_3_2_6 <= _GEN_9619;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_3_2_6 <= _GEN_5523; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_6 <= 1'h0;
      end else begin
        mask_3_2_6 <= _GEN_1379;
      end
    end else begin
      mask_3_2_6 <= _GEN_1379;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_3_2_7 <= _GEN_9683;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_3_2_7 <= _GEN_5587; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_2_7 <= 1'h0;
      end else begin
        mask_3_2_7 <= _GEN_1395;
      end
    end else begin
      mask_3_2_7 <= _GEN_1395;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_3_3_0 <= _GEN_9747;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_3_3_0 <= _GEN_5651; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_0 <= 1'h0;
      end else begin
        mask_3_3_0 <= _GEN_1411;
      end
    end else begin
      mask_3_3_0 <= _GEN_1411;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_3_3_1 <= _GEN_9811;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_3_3_1 <= _GEN_5715; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_1 <= 1'h0;
      end else begin
        mask_3_3_1 <= _GEN_1427;
      end
    end else begin
      mask_3_3_1 <= _GEN_1427;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_3_3_2 <= _GEN_9875;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_3_3_2 <= _GEN_5779; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_2 <= 1'h0;
      end else begin
        mask_3_3_2 <= _GEN_1443;
      end
    end else begin
      mask_3_3_2 <= _GEN_1443;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_3_3_3 <= _GEN_9939;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_3_3_3 <= _GEN_5843; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_3 <= 1'h0;
      end else begin
        mask_3_3_3 <= _GEN_1459;
      end
    end else begin
      mask_3_3_3 <= _GEN_1459;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_3_3_4 <= _GEN_10003;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_3_3_4 <= _GEN_5907; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_4 <= 1'h0;
      end else begin
        mask_3_3_4 <= _GEN_1475;
      end
    end else begin
      mask_3_3_4 <= _GEN_1475;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_3_3_5 <= _GEN_10067;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_3_3_5 <= _GEN_5971; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_5 <= 1'h0;
      end else begin
        mask_3_3_5 <= _GEN_1491;
      end
    end else begin
      mask_3_3_5 <= _GEN_1491;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_3_3_6 <= _GEN_10131;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_3_3_6 <= _GEN_6035; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_6 <= 1'h0;
      end else begin
        mask_3_3_6 <= _GEN_1507;
      end
    end else begin
      mask_3_3_6 <= _GEN_1507;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_3_3_7 <= _GEN_10195;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_3_3_7 <= _GEN_6099; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_3_7 <= 1'h0;
      end else begin
        mask_3_3_7 <= _GEN_1523;
      end
    end else begin
      mask_3_3_7 <= _GEN_1523;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_3_4_0 <= _GEN_10259;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_3_4_0 <= _GEN_6163; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_0 <= 1'h0;
      end else begin
        mask_3_4_0 <= _GEN_1539;
      end
    end else begin
      mask_3_4_0 <= _GEN_1539;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_3_4_1 <= _GEN_10323;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_3_4_1 <= _GEN_6227; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_1 <= 1'h0;
      end else begin
        mask_3_4_1 <= _GEN_1555;
      end
    end else begin
      mask_3_4_1 <= _GEN_1555;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_3_4_2 <= _GEN_10387;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_3_4_2 <= _GEN_6291; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_2 <= 1'h0;
      end else begin
        mask_3_4_2 <= _GEN_1571;
      end
    end else begin
      mask_3_4_2 <= _GEN_1571;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_3_4_3 <= _GEN_10451;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_3_4_3 <= _GEN_6355; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_3 <= 1'h0;
      end else begin
        mask_3_4_3 <= _GEN_1587;
      end
    end else begin
      mask_3_4_3 <= _GEN_1587;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_3_4_4 <= _GEN_10515;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_3_4_4 <= _GEN_6419; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_4 <= 1'h0;
      end else begin
        mask_3_4_4 <= _GEN_1603;
      end
    end else begin
      mask_3_4_4 <= _GEN_1603;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_3_4_5 <= _GEN_10579;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_3_4_5 <= _GEN_6483; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_5 <= 1'h0;
      end else begin
        mask_3_4_5 <= _GEN_1619;
      end
    end else begin
      mask_3_4_5 <= _GEN_1619;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_3_4_6 <= _GEN_10643;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_3_4_6 <= _GEN_6547; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_6 <= 1'h0;
      end else begin
        mask_3_4_6 <= _GEN_1635;
      end
    end else begin
      mask_3_4_6 <= _GEN_1635;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_3_4_7 <= _GEN_10707;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_3_4_7 <= _GEN_6611; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_4_7 <= 1'h0;
      end else begin
        mask_3_4_7 <= _GEN_1651;
      end
    end else begin
      mask_3_4_7 <= _GEN_1651;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_3_5_0 <= _GEN_10771;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_3_5_0 <= _GEN_6675; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_0 <= 1'h0;
      end else begin
        mask_3_5_0 <= _GEN_1667;
      end
    end else begin
      mask_3_5_0 <= _GEN_1667;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_3_5_1 <= _GEN_10835;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_3_5_1 <= _GEN_6739; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_1 <= 1'h0;
      end else begin
        mask_3_5_1 <= _GEN_1683;
      end
    end else begin
      mask_3_5_1 <= _GEN_1683;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_3_5_2 <= _GEN_10899;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_3_5_2 <= _GEN_6803; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_2 <= 1'h0;
      end else begin
        mask_3_5_2 <= _GEN_1699;
      end
    end else begin
      mask_3_5_2 <= _GEN_1699;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_3_5_3 <= _GEN_10963;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_3_5_3 <= _GEN_6867; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_3 <= 1'h0;
      end else begin
        mask_3_5_3 <= _GEN_1715;
      end
    end else begin
      mask_3_5_3 <= _GEN_1715;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_3_5_4 <= _GEN_11027;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_3_5_4 <= _GEN_6931; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_4 <= 1'h0;
      end else begin
        mask_3_5_4 <= _GEN_1731;
      end
    end else begin
      mask_3_5_4 <= _GEN_1731;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_3_5_5 <= _GEN_11091;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_3_5_5 <= _GEN_6995; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_5 <= 1'h0;
      end else begin
        mask_3_5_5 <= _GEN_1747;
      end
    end else begin
      mask_3_5_5 <= _GEN_1747;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_3_5_6 <= _GEN_11155;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_3_5_6 <= _GEN_7059; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_6 <= 1'h0;
      end else begin
        mask_3_5_6 <= _GEN_1763;
      end
    end else begin
      mask_3_5_6 <= _GEN_1763;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_3_5_7 <= _GEN_11219;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_3_5_7 <= _GEN_7123; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_5_7 <= 1'h0;
      end else begin
        mask_3_5_7 <= _GEN_1779;
      end
    end else begin
      mask_3_5_7 <= _GEN_1779;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_3_6_0 <= _GEN_11283;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_3_6_0 <= _GEN_7187; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_0 <= 1'h0;
      end else begin
        mask_3_6_0 <= _GEN_1795;
      end
    end else begin
      mask_3_6_0 <= _GEN_1795;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_3_6_1 <= _GEN_11347;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_3_6_1 <= _GEN_7251; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_1 <= 1'h0;
      end else begin
        mask_3_6_1 <= _GEN_1811;
      end
    end else begin
      mask_3_6_1 <= _GEN_1811;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_3_6_2 <= _GEN_11411;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_3_6_2 <= _GEN_7315; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_2 <= 1'h0;
      end else begin
        mask_3_6_2 <= _GEN_1827;
      end
    end else begin
      mask_3_6_2 <= _GEN_1827;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_3_6_3 <= _GEN_11475;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_3_6_3 <= _GEN_7379; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_3 <= 1'h0;
      end else begin
        mask_3_6_3 <= _GEN_1843;
      end
    end else begin
      mask_3_6_3 <= _GEN_1843;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_3_6_4 <= _GEN_11539;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_3_6_4 <= _GEN_7443; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_4 <= 1'h0;
      end else begin
        mask_3_6_4 <= _GEN_1859;
      end
    end else begin
      mask_3_6_4 <= _GEN_1859;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_3_6_5 <= _GEN_11603;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_3_6_5 <= _GEN_7507; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_5 <= 1'h0;
      end else begin
        mask_3_6_5 <= _GEN_1875;
      end
    end else begin
      mask_3_6_5 <= _GEN_1875;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_3_6_6 <= _GEN_11667;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_3_6_6 <= _GEN_7571; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_6 <= 1'h0;
      end else begin
        mask_3_6_6 <= _GEN_1891;
      end
    end else begin
      mask_3_6_6 <= _GEN_1891;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_3_6_7 <= _GEN_11731;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_3_6_7 <= _GEN_7635; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_6_7 <= 1'h0;
      end else begin
        mask_3_6_7 <= _GEN_1907;
      end
    end else begin
      mask_3_6_7 <= _GEN_1907;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_3_7_0 <= _GEN_11795;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_3_7_0 <= _GEN_7699; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_0 <= 1'h0;
      end else begin
        mask_3_7_0 <= _GEN_1923;
      end
    end else begin
      mask_3_7_0 <= _GEN_1923;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_3_7_1 <= _GEN_11859;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_3_7_1 <= _GEN_7763; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_1 <= 1'h0;
      end else begin
        mask_3_7_1 <= _GEN_1939;
      end
    end else begin
      mask_3_7_1 <= _GEN_1939;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_3_7_2 <= _GEN_11923;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_3_7_2 <= _GEN_7827; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_2 <= 1'h0;
      end else begin
        mask_3_7_2 <= _GEN_1955;
      end
    end else begin
      mask_3_7_2 <= _GEN_1955;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_3_7_3 <= _GEN_11987;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_3_7_3 <= _GEN_7891; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_3 <= 1'h0;
      end else begin
        mask_3_7_3 <= _GEN_1971;
      end
    end else begin
      mask_3_7_3 <= _GEN_1971;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_3_7_4 <= _GEN_12051;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_3_7_4 <= _GEN_7955; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_4 <= 1'h0;
      end else begin
        mask_3_7_4 <= _GEN_1987;
      end
    end else begin
      mask_3_7_4 <= _GEN_1987;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_3_7_5 <= _GEN_12115;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_3_7_5 <= _GEN_8019; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_5 <= 1'h0;
      end else begin
        mask_3_7_5 <= _GEN_2003;
      end
    end else begin
      mask_3_7_5 <= _GEN_2003;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_3_7_6 <= _GEN_12179;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_3_7_6 <= _GEN_8083; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_6 <= 1'h0;
      end else begin
        mask_3_7_6 <= _GEN_2019;
      end
    end else begin
      mask_3_7_6 <= _GEN_2019;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_3_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_3_7_7 <= _GEN_12243;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_3_7_7 <= _GEN_8147; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h3 == line_mask_clean_line_1) begin
        mask_3_7_7 <= 1'h0;
      end else begin
        mask_3_7_7 <= _GEN_2035;
      end
    end else begin
      mask_3_7_7 <= _GEN_2035;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_4_0_0 <= _GEN_8212;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_4_0_0 <= _GEN_4116; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_0 <= 1'h0;
      end else begin
        mask_4_0_0 <= _GEN_1028;
      end
    end else begin
      mask_4_0_0 <= _GEN_1028;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_4_0_1 <= _GEN_8276;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_4_0_1 <= _GEN_4180; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_1 <= 1'h0;
      end else begin
        mask_4_0_1 <= _GEN_1044;
      end
    end else begin
      mask_4_0_1 <= _GEN_1044;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_4_0_2 <= _GEN_8340;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_4_0_2 <= _GEN_4244; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_2 <= 1'h0;
      end else begin
        mask_4_0_2 <= _GEN_1060;
      end
    end else begin
      mask_4_0_2 <= _GEN_1060;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_4_0_3 <= _GEN_8404;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_4_0_3 <= _GEN_4308; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_3 <= 1'h0;
      end else begin
        mask_4_0_3 <= _GEN_1076;
      end
    end else begin
      mask_4_0_3 <= _GEN_1076;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_4_0_4 <= _GEN_8468;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_4_0_4 <= _GEN_4372; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_4 <= 1'h0;
      end else begin
        mask_4_0_4 <= _GEN_1092;
      end
    end else begin
      mask_4_0_4 <= _GEN_1092;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_4_0_5 <= _GEN_8532;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_4_0_5 <= _GEN_4436; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_5 <= 1'h0;
      end else begin
        mask_4_0_5 <= _GEN_1108;
      end
    end else begin
      mask_4_0_5 <= _GEN_1108;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_4_0_6 <= _GEN_8596;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_4_0_6 <= _GEN_4500; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_6 <= 1'h0;
      end else begin
        mask_4_0_6 <= _GEN_1124;
      end
    end else begin
      mask_4_0_6 <= _GEN_1124;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_4_0_7 <= _GEN_8660;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_4_0_7 <= _GEN_4564; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_0_7 <= 1'h0;
      end else begin
        mask_4_0_7 <= _GEN_1140;
      end
    end else begin
      mask_4_0_7 <= _GEN_1140;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_4_1_0 <= _GEN_8724;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_4_1_0 <= _GEN_4628; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_0 <= 1'h0;
      end else begin
        mask_4_1_0 <= _GEN_1156;
      end
    end else begin
      mask_4_1_0 <= _GEN_1156;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_4_1_1 <= _GEN_8788;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_4_1_1 <= _GEN_4692; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_1 <= 1'h0;
      end else begin
        mask_4_1_1 <= _GEN_1172;
      end
    end else begin
      mask_4_1_1 <= _GEN_1172;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_4_1_2 <= _GEN_8852;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_4_1_2 <= _GEN_4756; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_2 <= 1'h0;
      end else begin
        mask_4_1_2 <= _GEN_1188;
      end
    end else begin
      mask_4_1_2 <= _GEN_1188;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_4_1_3 <= _GEN_8916;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_4_1_3 <= _GEN_4820; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_3 <= 1'h0;
      end else begin
        mask_4_1_3 <= _GEN_1204;
      end
    end else begin
      mask_4_1_3 <= _GEN_1204;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_4_1_4 <= _GEN_8980;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_4_1_4 <= _GEN_4884; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_4 <= 1'h0;
      end else begin
        mask_4_1_4 <= _GEN_1220;
      end
    end else begin
      mask_4_1_4 <= _GEN_1220;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_4_1_5 <= _GEN_9044;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_4_1_5 <= _GEN_4948; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_5 <= 1'h0;
      end else begin
        mask_4_1_5 <= _GEN_1236;
      end
    end else begin
      mask_4_1_5 <= _GEN_1236;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_4_1_6 <= _GEN_9108;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_4_1_6 <= _GEN_5012; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_6 <= 1'h0;
      end else begin
        mask_4_1_6 <= _GEN_1252;
      end
    end else begin
      mask_4_1_6 <= _GEN_1252;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_4_1_7 <= _GEN_9172;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_4_1_7 <= _GEN_5076; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_1_7 <= 1'h0;
      end else begin
        mask_4_1_7 <= _GEN_1268;
      end
    end else begin
      mask_4_1_7 <= _GEN_1268;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_4_2_0 <= _GEN_9236;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_4_2_0 <= _GEN_5140; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_0 <= 1'h0;
      end else begin
        mask_4_2_0 <= _GEN_1284;
      end
    end else begin
      mask_4_2_0 <= _GEN_1284;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_4_2_1 <= _GEN_9300;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_4_2_1 <= _GEN_5204; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_1 <= 1'h0;
      end else begin
        mask_4_2_1 <= _GEN_1300;
      end
    end else begin
      mask_4_2_1 <= _GEN_1300;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_4_2_2 <= _GEN_9364;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_4_2_2 <= _GEN_5268; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_2 <= 1'h0;
      end else begin
        mask_4_2_2 <= _GEN_1316;
      end
    end else begin
      mask_4_2_2 <= _GEN_1316;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_4_2_3 <= _GEN_9428;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_4_2_3 <= _GEN_5332; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_3 <= 1'h0;
      end else begin
        mask_4_2_3 <= _GEN_1332;
      end
    end else begin
      mask_4_2_3 <= _GEN_1332;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_4_2_4 <= _GEN_9492;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_4_2_4 <= _GEN_5396; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_4 <= 1'h0;
      end else begin
        mask_4_2_4 <= _GEN_1348;
      end
    end else begin
      mask_4_2_4 <= _GEN_1348;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_4_2_5 <= _GEN_9556;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_4_2_5 <= _GEN_5460; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_5 <= 1'h0;
      end else begin
        mask_4_2_5 <= _GEN_1364;
      end
    end else begin
      mask_4_2_5 <= _GEN_1364;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_4_2_6 <= _GEN_9620;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_4_2_6 <= _GEN_5524; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_6 <= 1'h0;
      end else begin
        mask_4_2_6 <= _GEN_1380;
      end
    end else begin
      mask_4_2_6 <= _GEN_1380;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_4_2_7 <= _GEN_9684;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_4_2_7 <= _GEN_5588; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_2_7 <= 1'h0;
      end else begin
        mask_4_2_7 <= _GEN_1396;
      end
    end else begin
      mask_4_2_7 <= _GEN_1396;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_4_3_0 <= _GEN_9748;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_4_3_0 <= _GEN_5652; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_0 <= 1'h0;
      end else begin
        mask_4_3_0 <= _GEN_1412;
      end
    end else begin
      mask_4_3_0 <= _GEN_1412;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_4_3_1 <= _GEN_9812;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_4_3_1 <= _GEN_5716; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_1 <= 1'h0;
      end else begin
        mask_4_3_1 <= _GEN_1428;
      end
    end else begin
      mask_4_3_1 <= _GEN_1428;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_4_3_2 <= _GEN_9876;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_4_3_2 <= _GEN_5780; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_2 <= 1'h0;
      end else begin
        mask_4_3_2 <= _GEN_1444;
      end
    end else begin
      mask_4_3_2 <= _GEN_1444;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_4_3_3 <= _GEN_9940;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_4_3_3 <= _GEN_5844; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_3 <= 1'h0;
      end else begin
        mask_4_3_3 <= _GEN_1460;
      end
    end else begin
      mask_4_3_3 <= _GEN_1460;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_4_3_4 <= _GEN_10004;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_4_3_4 <= _GEN_5908; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_4 <= 1'h0;
      end else begin
        mask_4_3_4 <= _GEN_1476;
      end
    end else begin
      mask_4_3_4 <= _GEN_1476;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_4_3_5 <= _GEN_10068;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_4_3_5 <= _GEN_5972; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_5 <= 1'h0;
      end else begin
        mask_4_3_5 <= _GEN_1492;
      end
    end else begin
      mask_4_3_5 <= _GEN_1492;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_4_3_6 <= _GEN_10132;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_4_3_6 <= _GEN_6036; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_6 <= 1'h0;
      end else begin
        mask_4_3_6 <= _GEN_1508;
      end
    end else begin
      mask_4_3_6 <= _GEN_1508;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_4_3_7 <= _GEN_10196;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_4_3_7 <= _GEN_6100; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_3_7 <= 1'h0;
      end else begin
        mask_4_3_7 <= _GEN_1524;
      end
    end else begin
      mask_4_3_7 <= _GEN_1524;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_4_4_0 <= _GEN_10260;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_4_4_0 <= _GEN_6164; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_0 <= 1'h0;
      end else begin
        mask_4_4_0 <= _GEN_1540;
      end
    end else begin
      mask_4_4_0 <= _GEN_1540;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_4_4_1 <= _GEN_10324;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_4_4_1 <= _GEN_6228; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_1 <= 1'h0;
      end else begin
        mask_4_4_1 <= _GEN_1556;
      end
    end else begin
      mask_4_4_1 <= _GEN_1556;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_4_4_2 <= _GEN_10388;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_4_4_2 <= _GEN_6292; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_2 <= 1'h0;
      end else begin
        mask_4_4_2 <= _GEN_1572;
      end
    end else begin
      mask_4_4_2 <= _GEN_1572;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_4_4_3 <= _GEN_10452;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_4_4_3 <= _GEN_6356; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_3 <= 1'h0;
      end else begin
        mask_4_4_3 <= _GEN_1588;
      end
    end else begin
      mask_4_4_3 <= _GEN_1588;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_4_4_4 <= _GEN_10516;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_4_4_4 <= _GEN_6420; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_4 <= 1'h0;
      end else begin
        mask_4_4_4 <= _GEN_1604;
      end
    end else begin
      mask_4_4_4 <= _GEN_1604;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_4_4_5 <= _GEN_10580;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_4_4_5 <= _GEN_6484; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_5 <= 1'h0;
      end else begin
        mask_4_4_5 <= _GEN_1620;
      end
    end else begin
      mask_4_4_5 <= _GEN_1620;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_4_4_6 <= _GEN_10644;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_4_4_6 <= _GEN_6548; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_6 <= 1'h0;
      end else begin
        mask_4_4_6 <= _GEN_1636;
      end
    end else begin
      mask_4_4_6 <= _GEN_1636;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_4_4_7 <= _GEN_10708;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_4_4_7 <= _GEN_6612; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_4_7 <= 1'h0;
      end else begin
        mask_4_4_7 <= _GEN_1652;
      end
    end else begin
      mask_4_4_7 <= _GEN_1652;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_4_5_0 <= _GEN_10772;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_4_5_0 <= _GEN_6676; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_0 <= 1'h0;
      end else begin
        mask_4_5_0 <= _GEN_1668;
      end
    end else begin
      mask_4_5_0 <= _GEN_1668;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_4_5_1 <= _GEN_10836;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_4_5_1 <= _GEN_6740; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_1 <= 1'h0;
      end else begin
        mask_4_5_1 <= _GEN_1684;
      end
    end else begin
      mask_4_5_1 <= _GEN_1684;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_4_5_2 <= _GEN_10900;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_4_5_2 <= _GEN_6804; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_2 <= 1'h0;
      end else begin
        mask_4_5_2 <= _GEN_1700;
      end
    end else begin
      mask_4_5_2 <= _GEN_1700;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_4_5_3 <= _GEN_10964;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_4_5_3 <= _GEN_6868; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_3 <= 1'h0;
      end else begin
        mask_4_5_3 <= _GEN_1716;
      end
    end else begin
      mask_4_5_3 <= _GEN_1716;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_4_5_4 <= _GEN_11028;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_4_5_4 <= _GEN_6932; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_4 <= 1'h0;
      end else begin
        mask_4_5_4 <= _GEN_1732;
      end
    end else begin
      mask_4_5_4 <= _GEN_1732;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_4_5_5 <= _GEN_11092;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_4_5_5 <= _GEN_6996; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_5 <= 1'h0;
      end else begin
        mask_4_5_5 <= _GEN_1748;
      end
    end else begin
      mask_4_5_5 <= _GEN_1748;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_4_5_6 <= _GEN_11156;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_4_5_6 <= _GEN_7060; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_6 <= 1'h0;
      end else begin
        mask_4_5_6 <= _GEN_1764;
      end
    end else begin
      mask_4_5_6 <= _GEN_1764;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_4_5_7 <= _GEN_11220;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_4_5_7 <= _GEN_7124; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_5_7 <= 1'h0;
      end else begin
        mask_4_5_7 <= _GEN_1780;
      end
    end else begin
      mask_4_5_7 <= _GEN_1780;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_4_6_0 <= _GEN_11284;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_4_6_0 <= _GEN_7188; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_0 <= 1'h0;
      end else begin
        mask_4_6_0 <= _GEN_1796;
      end
    end else begin
      mask_4_6_0 <= _GEN_1796;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_4_6_1 <= _GEN_11348;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_4_6_1 <= _GEN_7252; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_1 <= 1'h0;
      end else begin
        mask_4_6_1 <= _GEN_1812;
      end
    end else begin
      mask_4_6_1 <= _GEN_1812;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_4_6_2 <= _GEN_11412;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_4_6_2 <= _GEN_7316; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_2 <= 1'h0;
      end else begin
        mask_4_6_2 <= _GEN_1828;
      end
    end else begin
      mask_4_6_2 <= _GEN_1828;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_4_6_3 <= _GEN_11476;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_4_6_3 <= _GEN_7380; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_3 <= 1'h0;
      end else begin
        mask_4_6_3 <= _GEN_1844;
      end
    end else begin
      mask_4_6_3 <= _GEN_1844;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_4_6_4 <= _GEN_11540;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_4_6_4 <= _GEN_7444; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_4 <= 1'h0;
      end else begin
        mask_4_6_4 <= _GEN_1860;
      end
    end else begin
      mask_4_6_4 <= _GEN_1860;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_4_6_5 <= _GEN_11604;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_4_6_5 <= _GEN_7508; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_5 <= 1'h0;
      end else begin
        mask_4_6_5 <= _GEN_1876;
      end
    end else begin
      mask_4_6_5 <= _GEN_1876;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_4_6_6 <= _GEN_11668;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_4_6_6 <= _GEN_7572; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_6 <= 1'h0;
      end else begin
        mask_4_6_6 <= _GEN_1892;
      end
    end else begin
      mask_4_6_6 <= _GEN_1892;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_4_6_7 <= _GEN_11732;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_4_6_7 <= _GEN_7636; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_6_7 <= 1'h0;
      end else begin
        mask_4_6_7 <= _GEN_1908;
      end
    end else begin
      mask_4_6_7 <= _GEN_1908;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_4_7_0 <= _GEN_11796;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_4_7_0 <= _GEN_7700; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_0 <= 1'h0;
      end else begin
        mask_4_7_0 <= _GEN_1924;
      end
    end else begin
      mask_4_7_0 <= _GEN_1924;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_4_7_1 <= _GEN_11860;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_4_7_1 <= _GEN_7764; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_1 <= 1'h0;
      end else begin
        mask_4_7_1 <= _GEN_1940;
      end
    end else begin
      mask_4_7_1 <= _GEN_1940;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_4_7_2 <= _GEN_11924;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_4_7_2 <= _GEN_7828; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_2 <= 1'h0;
      end else begin
        mask_4_7_2 <= _GEN_1956;
      end
    end else begin
      mask_4_7_2 <= _GEN_1956;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_4_7_3 <= _GEN_11988;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_4_7_3 <= _GEN_7892; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_3 <= 1'h0;
      end else begin
        mask_4_7_3 <= _GEN_1972;
      end
    end else begin
      mask_4_7_3 <= _GEN_1972;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_4_7_4 <= _GEN_12052;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_4_7_4 <= _GEN_7956; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_4 <= 1'h0;
      end else begin
        mask_4_7_4 <= _GEN_1988;
      end
    end else begin
      mask_4_7_4 <= _GEN_1988;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_4_7_5 <= _GEN_12116;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_4_7_5 <= _GEN_8020; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_5 <= 1'h0;
      end else begin
        mask_4_7_5 <= _GEN_2004;
      end
    end else begin
      mask_4_7_5 <= _GEN_2004;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_4_7_6 <= _GEN_12180;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_4_7_6 <= _GEN_8084; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_6 <= 1'h0;
      end else begin
        mask_4_7_6 <= _GEN_2020;
      end
    end else begin
      mask_4_7_6 <= _GEN_2020;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_4_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_4_7_7 <= _GEN_12244;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_4_7_7 <= _GEN_8148; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h4 == line_mask_clean_line_1) begin
        mask_4_7_7 <= 1'h0;
      end else begin
        mask_4_7_7 <= _GEN_2036;
      end
    end else begin
      mask_4_7_7 <= _GEN_2036;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_5_0_0 <= _GEN_8213;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_5_0_0 <= _GEN_4117; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_0 <= 1'h0;
      end else begin
        mask_5_0_0 <= _GEN_1029;
      end
    end else begin
      mask_5_0_0 <= _GEN_1029;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_5_0_1 <= _GEN_8277;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_5_0_1 <= _GEN_4181; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_1 <= 1'h0;
      end else begin
        mask_5_0_1 <= _GEN_1045;
      end
    end else begin
      mask_5_0_1 <= _GEN_1045;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_5_0_2 <= _GEN_8341;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_5_0_2 <= _GEN_4245; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_2 <= 1'h0;
      end else begin
        mask_5_0_2 <= _GEN_1061;
      end
    end else begin
      mask_5_0_2 <= _GEN_1061;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_5_0_3 <= _GEN_8405;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_5_0_3 <= _GEN_4309; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_3 <= 1'h0;
      end else begin
        mask_5_0_3 <= _GEN_1077;
      end
    end else begin
      mask_5_0_3 <= _GEN_1077;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_5_0_4 <= _GEN_8469;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_5_0_4 <= _GEN_4373; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_4 <= 1'h0;
      end else begin
        mask_5_0_4 <= _GEN_1093;
      end
    end else begin
      mask_5_0_4 <= _GEN_1093;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_5_0_5 <= _GEN_8533;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_5_0_5 <= _GEN_4437; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_5 <= 1'h0;
      end else begin
        mask_5_0_5 <= _GEN_1109;
      end
    end else begin
      mask_5_0_5 <= _GEN_1109;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_5_0_6 <= _GEN_8597;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_5_0_6 <= _GEN_4501; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_6 <= 1'h0;
      end else begin
        mask_5_0_6 <= _GEN_1125;
      end
    end else begin
      mask_5_0_6 <= _GEN_1125;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_5_0_7 <= _GEN_8661;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_5_0_7 <= _GEN_4565; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_0_7 <= 1'h0;
      end else begin
        mask_5_0_7 <= _GEN_1141;
      end
    end else begin
      mask_5_0_7 <= _GEN_1141;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_5_1_0 <= _GEN_8725;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_5_1_0 <= _GEN_4629; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_0 <= 1'h0;
      end else begin
        mask_5_1_0 <= _GEN_1157;
      end
    end else begin
      mask_5_1_0 <= _GEN_1157;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_5_1_1 <= _GEN_8789;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_5_1_1 <= _GEN_4693; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_1 <= 1'h0;
      end else begin
        mask_5_1_1 <= _GEN_1173;
      end
    end else begin
      mask_5_1_1 <= _GEN_1173;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_5_1_2 <= _GEN_8853;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_5_1_2 <= _GEN_4757; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_2 <= 1'h0;
      end else begin
        mask_5_1_2 <= _GEN_1189;
      end
    end else begin
      mask_5_1_2 <= _GEN_1189;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_5_1_3 <= _GEN_8917;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_5_1_3 <= _GEN_4821; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_3 <= 1'h0;
      end else begin
        mask_5_1_3 <= _GEN_1205;
      end
    end else begin
      mask_5_1_3 <= _GEN_1205;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_5_1_4 <= _GEN_8981;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_5_1_4 <= _GEN_4885; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_4 <= 1'h0;
      end else begin
        mask_5_1_4 <= _GEN_1221;
      end
    end else begin
      mask_5_1_4 <= _GEN_1221;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_5_1_5 <= _GEN_9045;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_5_1_5 <= _GEN_4949; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_5 <= 1'h0;
      end else begin
        mask_5_1_5 <= _GEN_1237;
      end
    end else begin
      mask_5_1_5 <= _GEN_1237;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_5_1_6 <= _GEN_9109;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_5_1_6 <= _GEN_5013; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_6 <= 1'h0;
      end else begin
        mask_5_1_6 <= _GEN_1253;
      end
    end else begin
      mask_5_1_6 <= _GEN_1253;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_5_1_7 <= _GEN_9173;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_5_1_7 <= _GEN_5077; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_1_7 <= 1'h0;
      end else begin
        mask_5_1_7 <= _GEN_1269;
      end
    end else begin
      mask_5_1_7 <= _GEN_1269;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_5_2_0 <= _GEN_9237;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_5_2_0 <= _GEN_5141; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_0 <= 1'h0;
      end else begin
        mask_5_2_0 <= _GEN_1285;
      end
    end else begin
      mask_5_2_0 <= _GEN_1285;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_5_2_1 <= _GEN_9301;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_5_2_1 <= _GEN_5205; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_1 <= 1'h0;
      end else begin
        mask_5_2_1 <= _GEN_1301;
      end
    end else begin
      mask_5_2_1 <= _GEN_1301;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_5_2_2 <= _GEN_9365;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_5_2_2 <= _GEN_5269; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_2 <= 1'h0;
      end else begin
        mask_5_2_2 <= _GEN_1317;
      end
    end else begin
      mask_5_2_2 <= _GEN_1317;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_5_2_3 <= _GEN_9429;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_5_2_3 <= _GEN_5333; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_3 <= 1'h0;
      end else begin
        mask_5_2_3 <= _GEN_1333;
      end
    end else begin
      mask_5_2_3 <= _GEN_1333;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_5_2_4 <= _GEN_9493;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_5_2_4 <= _GEN_5397; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_4 <= 1'h0;
      end else begin
        mask_5_2_4 <= _GEN_1349;
      end
    end else begin
      mask_5_2_4 <= _GEN_1349;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_5_2_5 <= _GEN_9557;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_5_2_5 <= _GEN_5461; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_5 <= 1'h0;
      end else begin
        mask_5_2_5 <= _GEN_1365;
      end
    end else begin
      mask_5_2_5 <= _GEN_1365;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_5_2_6 <= _GEN_9621;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_5_2_6 <= _GEN_5525; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_6 <= 1'h0;
      end else begin
        mask_5_2_6 <= _GEN_1381;
      end
    end else begin
      mask_5_2_6 <= _GEN_1381;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_5_2_7 <= _GEN_9685;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_5_2_7 <= _GEN_5589; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_2_7 <= 1'h0;
      end else begin
        mask_5_2_7 <= _GEN_1397;
      end
    end else begin
      mask_5_2_7 <= _GEN_1397;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_5_3_0 <= _GEN_9749;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_5_3_0 <= _GEN_5653; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_0 <= 1'h0;
      end else begin
        mask_5_3_0 <= _GEN_1413;
      end
    end else begin
      mask_5_3_0 <= _GEN_1413;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_5_3_1 <= _GEN_9813;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_5_3_1 <= _GEN_5717; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_1 <= 1'h0;
      end else begin
        mask_5_3_1 <= _GEN_1429;
      end
    end else begin
      mask_5_3_1 <= _GEN_1429;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_5_3_2 <= _GEN_9877;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_5_3_2 <= _GEN_5781; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_2 <= 1'h0;
      end else begin
        mask_5_3_2 <= _GEN_1445;
      end
    end else begin
      mask_5_3_2 <= _GEN_1445;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_5_3_3 <= _GEN_9941;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_5_3_3 <= _GEN_5845; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_3 <= 1'h0;
      end else begin
        mask_5_3_3 <= _GEN_1461;
      end
    end else begin
      mask_5_3_3 <= _GEN_1461;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_5_3_4 <= _GEN_10005;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_5_3_4 <= _GEN_5909; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_4 <= 1'h0;
      end else begin
        mask_5_3_4 <= _GEN_1477;
      end
    end else begin
      mask_5_3_4 <= _GEN_1477;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_5_3_5 <= _GEN_10069;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_5_3_5 <= _GEN_5973; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_5 <= 1'h0;
      end else begin
        mask_5_3_5 <= _GEN_1493;
      end
    end else begin
      mask_5_3_5 <= _GEN_1493;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_5_3_6 <= _GEN_10133;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_5_3_6 <= _GEN_6037; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_6 <= 1'h0;
      end else begin
        mask_5_3_6 <= _GEN_1509;
      end
    end else begin
      mask_5_3_6 <= _GEN_1509;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_5_3_7 <= _GEN_10197;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_5_3_7 <= _GEN_6101; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_3_7 <= 1'h0;
      end else begin
        mask_5_3_7 <= _GEN_1525;
      end
    end else begin
      mask_5_3_7 <= _GEN_1525;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_5_4_0 <= _GEN_10261;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_5_4_0 <= _GEN_6165; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_0 <= 1'h0;
      end else begin
        mask_5_4_0 <= _GEN_1541;
      end
    end else begin
      mask_5_4_0 <= _GEN_1541;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_5_4_1 <= _GEN_10325;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_5_4_1 <= _GEN_6229; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_1 <= 1'h0;
      end else begin
        mask_5_4_1 <= _GEN_1557;
      end
    end else begin
      mask_5_4_1 <= _GEN_1557;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_5_4_2 <= _GEN_10389;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_5_4_2 <= _GEN_6293; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_2 <= 1'h0;
      end else begin
        mask_5_4_2 <= _GEN_1573;
      end
    end else begin
      mask_5_4_2 <= _GEN_1573;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_5_4_3 <= _GEN_10453;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_5_4_3 <= _GEN_6357; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_3 <= 1'h0;
      end else begin
        mask_5_4_3 <= _GEN_1589;
      end
    end else begin
      mask_5_4_3 <= _GEN_1589;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_5_4_4 <= _GEN_10517;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_5_4_4 <= _GEN_6421; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_4 <= 1'h0;
      end else begin
        mask_5_4_4 <= _GEN_1605;
      end
    end else begin
      mask_5_4_4 <= _GEN_1605;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_5_4_5 <= _GEN_10581;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_5_4_5 <= _GEN_6485; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_5 <= 1'h0;
      end else begin
        mask_5_4_5 <= _GEN_1621;
      end
    end else begin
      mask_5_4_5 <= _GEN_1621;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_5_4_6 <= _GEN_10645;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_5_4_6 <= _GEN_6549; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_6 <= 1'h0;
      end else begin
        mask_5_4_6 <= _GEN_1637;
      end
    end else begin
      mask_5_4_6 <= _GEN_1637;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_5_4_7 <= _GEN_10709;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_5_4_7 <= _GEN_6613; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_4_7 <= 1'h0;
      end else begin
        mask_5_4_7 <= _GEN_1653;
      end
    end else begin
      mask_5_4_7 <= _GEN_1653;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_5_5_0 <= _GEN_10773;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_5_5_0 <= _GEN_6677; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_0 <= 1'h0;
      end else begin
        mask_5_5_0 <= _GEN_1669;
      end
    end else begin
      mask_5_5_0 <= _GEN_1669;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_5_5_1 <= _GEN_10837;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_5_5_1 <= _GEN_6741; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_1 <= 1'h0;
      end else begin
        mask_5_5_1 <= _GEN_1685;
      end
    end else begin
      mask_5_5_1 <= _GEN_1685;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_5_5_2 <= _GEN_10901;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_5_5_2 <= _GEN_6805; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_2 <= 1'h0;
      end else begin
        mask_5_5_2 <= _GEN_1701;
      end
    end else begin
      mask_5_5_2 <= _GEN_1701;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_5_5_3 <= _GEN_10965;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_5_5_3 <= _GEN_6869; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_3 <= 1'h0;
      end else begin
        mask_5_5_3 <= _GEN_1717;
      end
    end else begin
      mask_5_5_3 <= _GEN_1717;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_5_5_4 <= _GEN_11029;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_5_5_4 <= _GEN_6933; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_4 <= 1'h0;
      end else begin
        mask_5_5_4 <= _GEN_1733;
      end
    end else begin
      mask_5_5_4 <= _GEN_1733;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_5_5_5 <= _GEN_11093;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_5_5_5 <= _GEN_6997; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_5 <= 1'h0;
      end else begin
        mask_5_5_5 <= _GEN_1749;
      end
    end else begin
      mask_5_5_5 <= _GEN_1749;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_5_5_6 <= _GEN_11157;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_5_5_6 <= _GEN_7061; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_6 <= 1'h0;
      end else begin
        mask_5_5_6 <= _GEN_1765;
      end
    end else begin
      mask_5_5_6 <= _GEN_1765;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_5_5_7 <= _GEN_11221;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_5_5_7 <= _GEN_7125; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_5_7 <= 1'h0;
      end else begin
        mask_5_5_7 <= _GEN_1781;
      end
    end else begin
      mask_5_5_7 <= _GEN_1781;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_5_6_0 <= _GEN_11285;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_5_6_0 <= _GEN_7189; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_0 <= 1'h0;
      end else begin
        mask_5_6_0 <= _GEN_1797;
      end
    end else begin
      mask_5_6_0 <= _GEN_1797;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_5_6_1 <= _GEN_11349;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_5_6_1 <= _GEN_7253; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_1 <= 1'h0;
      end else begin
        mask_5_6_1 <= _GEN_1813;
      end
    end else begin
      mask_5_6_1 <= _GEN_1813;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_5_6_2 <= _GEN_11413;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_5_6_2 <= _GEN_7317; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_2 <= 1'h0;
      end else begin
        mask_5_6_2 <= _GEN_1829;
      end
    end else begin
      mask_5_6_2 <= _GEN_1829;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_5_6_3 <= _GEN_11477;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_5_6_3 <= _GEN_7381; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_3 <= 1'h0;
      end else begin
        mask_5_6_3 <= _GEN_1845;
      end
    end else begin
      mask_5_6_3 <= _GEN_1845;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_5_6_4 <= _GEN_11541;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_5_6_4 <= _GEN_7445; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_4 <= 1'h0;
      end else begin
        mask_5_6_4 <= _GEN_1861;
      end
    end else begin
      mask_5_6_4 <= _GEN_1861;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_5_6_5 <= _GEN_11605;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_5_6_5 <= _GEN_7509; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_5 <= 1'h0;
      end else begin
        mask_5_6_5 <= _GEN_1877;
      end
    end else begin
      mask_5_6_5 <= _GEN_1877;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_5_6_6 <= _GEN_11669;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_5_6_6 <= _GEN_7573; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_6 <= 1'h0;
      end else begin
        mask_5_6_6 <= _GEN_1893;
      end
    end else begin
      mask_5_6_6 <= _GEN_1893;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_5_6_7 <= _GEN_11733;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_5_6_7 <= _GEN_7637; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_6_7 <= 1'h0;
      end else begin
        mask_5_6_7 <= _GEN_1909;
      end
    end else begin
      mask_5_6_7 <= _GEN_1909;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_5_7_0 <= _GEN_11797;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_5_7_0 <= _GEN_7701; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_0 <= 1'h0;
      end else begin
        mask_5_7_0 <= _GEN_1925;
      end
    end else begin
      mask_5_7_0 <= _GEN_1925;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_5_7_1 <= _GEN_11861;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_5_7_1 <= _GEN_7765; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_1 <= 1'h0;
      end else begin
        mask_5_7_1 <= _GEN_1941;
      end
    end else begin
      mask_5_7_1 <= _GEN_1941;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_5_7_2 <= _GEN_11925;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_5_7_2 <= _GEN_7829; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_2 <= 1'h0;
      end else begin
        mask_5_7_2 <= _GEN_1957;
      end
    end else begin
      mask_5_7_2 <= _GEN_1957;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_5_7_3 <= _GEN_11989;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_5_7_3 <= _GEN_7893; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_3 <= 1'h0;
      end else begin
        mask_5_7_3 <= _GEN_1973;
      end
    end else begin
      mask_5_7_3 <= _GEN_1973;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_5_7_4 <= _GEN_12053;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_5_7_4 <= _GEN_7957; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_4 <= 1'h0;
      end else begin
        mask_5_7_4 <= _GEN_1989;
      end
    end else begin
      mask_5_7_4 <= _GEN_1989;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_5_7_5 <= _GEN_12117;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_5_7_5 <= _GEN_8021; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_5 <= 1'h0;
      end else begin
        mask_5_7_5 <= _GEN_2005;
      end
    end else begin
      mask_5_7_5 <= _GEN_2005;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_5_7_6 <= _GEN_12181;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_5_7_6 <= _GEN_8085; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_6 <= 1'h0;
      end else begin
        mask_5_7_6 <= _GEN_2021;
      end
    end else begin
      mask_5_7_6 <= _GEN_2021;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_5_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_5_7_7 <= _GEN_12245;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_5_7_7 <= _GEN_8149; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h5 == line_mask_clean_line_1) begin
        mask_5_7_7 <= 1'h0;
      end else begin
        mask_5_7_7 <= _GEN_2037;
      end
    end else begin
      mask_5_7_7 <= _GEN_2037;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_6_0_0 <= _GEN_8214;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_6_0_0 <= _GEN_4118; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_0 <= 1'h0;
      end else begin
        mask_6_0_0 <= _GEN_1030;
      end
    end else begin
      mask_6_0_0 <= _GEN_1030;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_6_0_1 <= _GEN_8278;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_6_0_1 <= _GEN_4182; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_1 <= 1'h0;
      end else begin
        mask_6_0_1 <= _GEN_1046;
      end
    end else begin
      mask_6_0_1 <= _GEN_1046;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_6_0_2 <= _GEN_8342;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_6_0_2 <= _GEN_4246; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_2 <= 1'h0;
      end else begin
        mask_6_0_2 <= _GEN_1062;
      end
    end else begin
      mask_6_0_2 <= _GEN_1062;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_6_0_3 <= _GEN_8406;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_6_0_3 <= _GEN_4310; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_3 <= 1'h0;
      end else begin
        mask_6_0_3 <= _GEN_1078;
      end
    end else begin
      mask_6_0_3 <= _GEN_1078;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_6_0_4 <= _GEN_8470;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_6_0_4 <= _GEN_4374; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_4 <= 1'h0;
      end else begin
        mask_6_0_4 <= _GEN_1094;
      end
    end else begin
      mask_6_0_4 <= _GEN_1094;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_6_0_5 <= _GEN_8534;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_6_0_5 <= _GEN_4438; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_5 <= 1'h0;
      end else begin
        mask_6_0_5 <= _GEN_1110;
      end
    end else begin
      mask_6_0_5 <= _GEN_1110;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_6_0_6 <= _GEN_8598;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_6_0_6 <= _GEN_4502; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_6 <= 1'h0;
      end else begin
        mask_6_0_6 <= _GEN_1126;
      end
    end else begin
      mask_6_0_6 <= _GEN_1126;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_6_0_7 <= _GEN_8662;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_6_0_7 <= _GEN_4566; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_0_7 <= 1'h0;
      end else begin
        mask_6_0_7 <= _GEN_1142;
      end
    end else begin
      mask_6_0_7 <= _GEN_1142;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_6_1_0 <= _GEN_8726;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_6_1_0 <= _GEN_4630; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_0 <= 1'h0;
      end else begin
        mask_6_1_0 <= _GEN_1158;
      end
    end else begin
      mask_6_1_0 <= _GEN_1158;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_6_1_1 <= _GEN_8790;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_6_1_1 <= _GEN_4694; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_1 <= 1'h0;
      end else begin
        mask_6_1_1 <= _GEN_1174;
      end
    end else begin
      mask_6_1_1 <= _GEN_1174;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_6_1_2 <= _GEN_8854;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_6_1_2 <= _GEN_4758; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_2 <= 1'h0;
      end else begin
        mask_6_1_2 <= _GEN_1190;
      end
    end else begin
      mask_6_1_2 <= _GEN_1190;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_6_1_3 <= _GEN_8918;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_6_1_3 <= _GEN_4822; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_3 <= 1'h0;
      end else begin
        mask_6_1_3 <= _GEN_1206;
      end
    end else begin
      mask_6_1_3 <= _GEN_1206;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_6_1_4 <= _GEN_8982;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_6_1_4 <= _GEN_4886; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_4 <= 1'h0;
      end else begin
        mask_6_1_4 <= _GEN_1222;
      end
    end else begin
      mask_6_1_4 <= _GEN_1222;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_6_1_5 <= _GEN_9046;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_6_1_5 <= _GEN_4950; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_5 <= 1'h0;
      end else begin
        mask_6_1_5 <= _GEN_1238;
      end
    end else begin
      mask_6_1_5 <= _GEN_1238;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_6_1_6 <= _GEN_9110;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_6_1_6 <= _GEN_5014; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_6 <= 1'h0;
      end else begin
        mask_6_1_6 <= _GEN_1254;
      end
    end else begin
      mask_6_1_6 <= _GEN_1254;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_6_1_7 <= _GEN_9174;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_6_1_7 <= _GEN_5078; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_1_7 <= 1'h0;
      end else begin
        mask_6_1_7 <= _GEN_1270;
      end
    end else begin
      mask_6_1_7 <= _GEN_1270;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_6_2_0 <= _GEN_9238;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_6_2_0 <= _GEN_5142; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_0 <= 1'h0;
      end else begin
        mask_6_2_0 <= _GEN_1286;
      end
    end else begin
      mask_6_2_0 <= _GEN_1286;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_6_2_1 <= _GEN_9302;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_6_2_1 <= _GEN_5206; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_1 <= 1'h0;
      end else begin
        mask_6_2_1 <= _GEN_1302;
      end
    end else begin
      mask_6_2_1 <= _GEN_1302;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_6_2_2 <= _GEN_9366;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_6_2_2 <= _GEN_5270; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_2 <= 1'h0;
      end else begin
        mask_6_2_2 <= _GEN_1318;
      end
    end else begin
      mask_6_2_2 <= _GEN_1318;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_6_2_3 <= _GEN_9430;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_6_2_3 <= _GEN_5334; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_3 <= 1'h0;
      end else begin
        mask_6_2_3 <= _GEN_1334;
      end
    end else begin
      mask_6_2_3 <= _GEN_1334;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_6_2_4 <= _GEN_9494;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_6_2_4 <= _GEN_5398; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_4 <= 1'h0;
      end else begin
        mask_6_2_4 <= _GEN_1350;
      end
    end else begin
      mask_6_2_4 <= _GEN_1350;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_6_2_5 <= _GEN_9558;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_6_2_5 <= _GEN_5462; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_5 <= 1'h0;
      end else begin
        mask_6_2_5 <= _GEN_1366;
      end
    end else begin
      mask_6_2_5 <= _GEN_1366;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_6_2_6 <= _GEN_9622;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_6_2_6 <= _GEN_5526; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_6 <= 1'h0;
      end else begin
        mask_6_2_6 <= _GEN_1382;
      end
    end else begin
      mask_6_2_6 <= _GEN_1382;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_6_2_7 <= _GEN_9686;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_6_2_7 <= _GEN_5590; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_2_7 <= 1'h0;
      end else begin
        mask_6_2_7 <= _GEN_1398;
      end
    end else begin
      mask_6_2_7 <= _GEN_1398;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_6_3_0 <= _GEN_9750;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_6_3_0 <= _GEN_5654; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_0 <= 1'h0;
      end else begin
        mask_6_3_0 <= _GEN_1414;
      end
    end else begin
      mask_6_3_0 <= _GEN_1414;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_6_3_1 <= _GEN_9814;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_6_3_1 <= _GEN_5718; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_1 <= 1'h0;
      end else begin
        mask_6_3_1 <= _GEN_1430;
      end
    end else begin
      mask_6_3_1 <= _GEN_1430;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_6_3_2 <= _GEN_9878;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_6_3_2 <= _GEN_5782; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_2 <= 1'h0;
      end else begin
        mask_6_3_2 <= _GEN_1446;
      end
    end else begin
      mask_6_3_2 <= _GEN_1446;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_6_3_3 <= _GEN_9942;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_6_3_3 <= _GEN_5846; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_3 <= 1'h0;
      end else begin
        mask_6_3_3 <= _GEN_1462;
      end
    end else begin
      mask_6_3_3 <= _GEN_1462;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_6_3_4 <= _GEN_10006;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_6_3_4 <= _GEN_5910; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_4 <= 1'h0;
      end else begin
        mask_6_3_4 <= _GEN_1478;
      end
    end else begin
      mask_6_3_4 <= _GEN_1478;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_6_3_5 <= _GEN_10070;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_6_3_5 <= _GEN_5974; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_5 <= 1'h0;
      end else begin
        mask_6_3_5 <= _GEN_1494;
      end
    end else begin
      mask_6_3_5 <= _GEN_1494;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_6_3_6 <= _GEN_10134;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_6_3_6 <= _GEN_6038; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_6 <= 1'h0;
      end else begin
        mask_6_3_6 <= _GEN_1510;
      end
    end else begin
      mask_6_3_6 <= _GEN_1510;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_6_3_7 <= _GEN_10198;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_6_3_7 <= _GEN_6102; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_3_7 <= 1'h0;
      end else begin
        mask_6_3_7 <= _GEN_1526;
      end
    end else begin
      mask_6_3_7 <= _GEN_1526;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_6_4_0 <= _GEN_10262;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_6_4_0 <= _GEN_6166; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_0 <= 1'h0;
      end else begin
        mask_6_4_0 <= _GEN_1542;
      end
    end else begin
      mask_6_4_0 <= _GEN_1542;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_6_4_1 <= _GEN_10326;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_6_4_1 <= _GEN_6230; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_1 <= 1'h0;
      end else begin
        mask_6_4_1 <= _GEN_1558;
      end
    end else begin
      mask_6_4_1 <= _GEN_1558;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_6_4_2 <= _GEN_10390;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_6_4_2 <= _GEN_6294; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_2 <= 1'h0;
      end else begin
        mask_6_4_2 <= _GEN_1574;
      end
    end else begin
      mask_6_4_2 <= _GEN_1574;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_6_4_3 <= _GEN_10454;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_6_4_3 <= _GEN_6358; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_3 <= 1'h0;
      end else begin
        mask_6_4_3 <= _GEN_1590;
      end
    end else begin
      mask_6_4_3 <= _GEN_1590;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_6_4_4 <= _GEN_10518;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_6_4_4 <= _GEN_6422; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_4 <= 1'h0;
      end else begin
        mask_6_4_4 <= _GEN_1606;
      end
    end else begin
      mask_6_4_4 <= _GEN_1606;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_6_4_5 <= _GEN_10582;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_6_4_5 <= _GEN_6486; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_5 <= 1'h0;
      end else begin
        mask_6_4_5 <= _GEN_1622;
      end
    end else begin
      mask_6_4_5 <= _GEN_1622;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_6_4_6 <= _GEN_10646;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_6_4_6 <= _GEN_6550; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_6 <= 1'h0;
      end else begin
        mask_6_4_6 <= _GEN_1638;
      end
    end else begin
      mask_6_4_6 <= _GEN_1638;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_6_4_7 <= _GEN_10710;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_6_4_7 <= _GEN_6614; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_4_7 <= 1'h0;
      end else begin
        mask_6_4_7 <= _GEN_1654;
      end
    end else begin
      mask_6_4_7 <= _GEN_1654;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_6_5_0 <= _GEN_10774;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_6_5_0 <= _GEN_6678; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_0 <= 1'h0;
      end else begin
        mask_6_5_0 <= _GEN_1670;
      end
    end else begin
      mask_6_5_0 <= _GEN_1670;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_6_5_1 <= _GEN_10838;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_6_5_1 <= _GEN_6742; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_1 <= 1'h0;
      end else begin
        mask_6_5_1 <= _GEN_1686;
      end
    end else begin
      mask_6_5_1 <= _GEN_1686;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_6_5_2 <= _GEN_10902;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_6_5_2 <= _GEN_6806; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_2 <= 1'h0;
      end else begin
        mask_6_5_2 <= _GEN_1702;
      end
    end else begin
      mask_6_5_2 <= _GEN_1702;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_6_5_3 <= _GEN_10966;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_6_5_3 <= _GEN_6870; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_3 <= 1'h0;
      end else begin
        mask_6_5_3 <= _GEN_1718;
      end
    end else begin
      mask_6_5_3 <= _GEN_1718;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_6_5_4 <= _GEN_11030;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_6_5_4 <= _GEN_6934; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_4 <= 1'h0;
      end else begin
        mask_6_5_4 <= _GEN_1734;
      end
    end else begin
      mask_6_5_4 <= _GEN_1734;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_6_5_5 <= _GEN_11094;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_6_5_5 <= _GEN_6998; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_5 <= 1'h0;
      end else begin
        mask_6_5_5 <= _GEN_1750;
      end
    end else begin
      mask_6_5_5 <= _GEN_1750;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_6_5_6 <= _GEN_11158;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_6_5_6 <= _GEN_7062; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_6 <= 1'h0;
      end else begin
        mask_6_5_6 <= _GEN_1766;
      end
    end else begin
      mask_6_5_6 <= _GEN_1766;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_6_5_7 <= _GEN_11222;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_6_5_7 <= _GEN_7126; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_5_7 <= 1'h0;
      end else begin
        mask_6_5_7 <= _GEN_1782;
      end
    end else begin
      mask_6_5_7 <= _GEN_1782;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_6_6_0 <= _GEN_11286;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_6_6_0 <= _GEN_7190; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_0 <= 1'h0;
      end else begin
        mask_6_6_0 <= _GEN_1798;
      end
    end else begin
      mask_6_6_0 <= _GEN_1798;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_6_6_1 <= _GEN_11350;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_6_6_1 <= _GEN_7254; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_1 <= 1'h0;
      end else begin
        mask_6_6_1 <= _GEN_1814;
      end
    end else begin
      mask_6_6_1 <= _GEN_1814;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_6_6_2 <= _GEN_11414;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_6_6_2 <= _GEN_7318; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_2 <= 1'h0;
      end else begin
        mask_6_6_2 <= _GEN_1830;
      end
    end else begin
      mask_6_6_2 <= _GEN_1830;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_6_6_3 <= _GEN_11478;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_6_6_3 <= _GEN_7382; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_3 <= 1'h0;
      end else begin
        mask_6_6_3 <= _GEN_1846;
      end
    end else begin
      mask_6_6_3 <= _GEN_1846;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_6_6_4 <= _GEN_11542;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_6_6_4 <= _GEN_7446; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_4 <= 1'h0;
      end else begin
        mask_6_6_4 <= _GEN_1862;
      end
    end else begin
      mask_6_6_4 <= _GEN_1862;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_6_6_5 <= _GEN_11606;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_6_6_5 <= _GEN_7510; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_5 <= 1'h0;
      end else begin
        mask_6_6_5 <= _GEN_1878;
      end
    end else begin
      mask_6_6_5 <= _GEN_1878;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_6_6_6 <= _GEN_11670;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_6_6_6 <= _GEN_7574; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_6 <= 1'h0;
      end else begin
        mask_6_6_6 <= _GEN_1894;
      end
    end else begin
      mask_6_6_6 <= _GEN_1894;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_6_6_7 <= _GEN_11734;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_6_6_7 <= _GEN_7638; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_6_7 <= 1'h0;
      end else begin
        mask_6_6_7 <= _GEN_1910;
      end
    end else begin
      mask_6_6_7 <= _GEN_1910;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_6_7_0 <= _GEN_11798;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_6_7_0 <= _GEN_7702; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_0 <= 1'h0;
      end else begin
        mask_6_7_0 <= _GEN_1926;
      end
    end else begin
      mask_6_7_0 <= _GEN_1926;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_6_7_1 <= _GEN_11862;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_6_7_1 <= _GEN_7766; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_1 <= 1'h0;
      end else begin
        mask_6_7_1 <= _GEN_1942;
      end
    end else begin
      mask_6_7_1 <= _GEN_1942;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_6_7_2 <= _GEN_11926;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_6_7_2 <= _GEN_7830; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_2 <= 1'h0;
      end else begin
        mask_6_7_2 <= _GEN_1958;
      end
    end else begin
      mask_6_7_2 <= _GEN_1958;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_6_7_3 <= _GEN_11990;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_6_7_3 <= _GEN_7894; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_3 <= 1'h0;
      end else begin
        mask_6_7_3 <= _GEN_1974;
      end
    end else begin
      mask_6_7_3 <= _GEN_1974;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_6_7_4 <= _GEN_12054;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_6_7_4 <= _GEN_7958; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_4 <= 1'h0;
      end else begin
        mask_6_7_4 <= _GEN_1990;
      end
    end else begin
      mask_6_7_4 <= _GEN_1990;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_6_7_5 <= _GEN_12118;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_6_7_5 <= _GEN_8022; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_5 <= 1'h0;
      end else begin
        mask_6_7_5 <= _GEN_2006;
      end
    end else begin
      mask_6_7_5 <= _GEN_2006;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_6_7_6 <= _GEN_12182;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_6_7_6 <= _GEN_8086; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_6 <= 1'h0;
      end else begin
        mask_6_7_6 <= _GEN_2022;
      end
    end else begin
      mask_6_7_6 <= _GEN_2022;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_6_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_6_7_7 <= _GEN_12246;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_6_7_7 <= _GEN_8150; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h6 == line_mask_clean_line_1) begin
        mask_6_7_7 <= 1'h0;
      end else begin
        mask_6_7_7 <= _GEN_2038;
      end
    end else begin
      mask_6_7_7 <= _GEN_2038;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_7_0_0 <= _GEN_8215;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_7_0_0 <= _GEN_4119; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_0 <= 1'h0;
      end else begin
        mask_7_0_0 <= _GEN_1031;
      end
    end else begin
      mask_7_0_0 <= _GEN_1031;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_7_0_1 <= _GEN_8279;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_7_0_1 <= _GEN_4183; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_1 <= 1'h0;
      end else begin
        mask_7_0_1 <= _GEN_1047;
      end
    end else begin
      mask_7_0_1 <= _GEN_1047;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_7_0_2 <= _GEN_8343;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_7_0_2 <= _GEN_4247; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_2 <= 1'h0;
      end else begin
        mask_7_0_2 <= _GEN_1063;
      end
    end else begin
      mask_7_0_2 <= _GEN_1063;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_7_0_3 <= _GEN_8407;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_7_0_3 <= _GEN_4311; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_3 <= 1'h0;
      end else begin
        mask_7_0_3 <= _GEN_1079;
      end
    end else begin
      mask_7_0_3 <= _GEN_1079;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_7_0_4 <= _GEN_8471;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_7_0_4 <= _GEN_4375; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_4 <= 1'h0;
      end else begin
        mask_7_0_4 <= _GEN_1095;
      end
    end else begin
      mask_7_0_4 <= _GEN_1095;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_7_0_5 <= _GEN_8535;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_7_0_5 <= _GEN_4439; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_5 <= 1'h0;
      end else begin
        mask_7_0_5 <= _GEN_1111;
      end
    end else begin
      mask_7_0_5 <= _GEN_1111;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_7_0_6 <= _GEN_8599;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_7_0_6 <= _GEN_4503; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_6 <= 1'h0;
      end else begin
        mask_7_0_6 <= _GEN_1127;
      end
    end else begin
      mask_7_0_6 <= _GEN_1127;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_7_0_7 <= _GEN_8663;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_7_0_7 <= _GEN_4567; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_0_7 <= 1'h0;
      end else begin
        mask_7_0_7 <= _GEN_1143;
      end
    end else begin
      mask_7_0_7 <= _GEN_1143;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_7_1_0 <= _GEN_8727;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_7_1_0 <= _GEN_4631; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_0 <= 1'h0;
      end else begin
        mask_7_1_0 <= _GEN_1159;
      end
    end else begin
      mask_7_1_0 <= _GEN_1159;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_7_1_1 <= _GEN_8791;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_7_1_1 <= _GEN_4695; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_1 <= 1'h0;
      end else begin
        mask_7_1_1 <= _GEN_1175;
      end
    end else begin
      mask_7_1_1 <= _GEN_1175;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_7_1_2 <= _GEN_8855;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_7_1_2 <= _GEN_4759; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_2 <= 1'h0;
      end else begin
        mask_7_1_2 <= _GEN_1191;
      end
    end else begin
      mask_7_1_2 <= _GEN_1191;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_7_1_3 <= _GEN_8919;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_7_1_3 <= _GEN_4823; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_3 <= 1'h0;
      end else begin
        mask_7_1_3 <= _GEN_1207;
      end
    end else begin
      mask_7_1_3 <= _GEN_1207;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_7_1_4 <= _GEN_8983;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_7_1_4 <= _GEN_4887; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_4 <= 1'h0;
      end else begin
        mask_7_1_4 <= _GEN_1223;
      end
    end else begin
      mask_7_1_4 <= _GEN_1223;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_7_1_5 <= _GEN_9047;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_7_1_5 <= _GEN_4951; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_5 <= 1'h0;
      end else begin
        mask_7_1_5 <= _GEN_1239;
      end
    end else begin
      mask_7_1_5 <= _GEN_1239;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_7_1_6 <= _GEN_9111;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_7_1_6 <= _GEN_5015; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_6 <= 1'h0;
      end else begin
        mask_7_1_6 <= _GEN_1255;
      end
    end else begin
      mask_7_1_6 <= _GEN_1255;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_7_1_7 <= _GEN_9175;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_7_1_7 <= _GEN_5079; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_1_7 <= 1'h0;
      end else begin
        mask_7_1_7 <= _GEN_1271;
      end
    end else begin
      mask_7_1_7 <= _GEN_1271;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_7_2_0 <= _GEN_9239;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_7_2_0 <= _GEN_5143; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_0 <= 1'h0;
      end else begin
        mask_7_2_0 <= _GEN_1287;
      end
    end else begin
      mask_7_2_0 <= _GEN_1287;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_7_2_1 <= _GEN_9303;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_7_2_1 <= _GEN_5207; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_1 <= 1'h0;
      end else begin
        mask_7_2_1 <= _GEN_1303;
      end
    end else begin
      mask_7_2_1 <= _GEN_1303;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_7_2_2 <= _GEN_9367;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_7_2_2 <= _GEN_5271; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_2 <= 1'h0;
      end else begin
        mask_7_2_2 <= _GEN_1319;
      end
    end else begin
      mask_7_2_2 <= _GEN_1319;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_7_2_3 <= _GEN_9431;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_7_2_3 <= _GEN_5335; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_3 <= 1'h0;
      end else begin
        mask_7_2_3 <= _GEN_1335;
      end
    end else begin
      mask_7_2_3 <= _GEN_1335;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_7_2_4 <= _GEN_9495;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_7_2_4 <= _GEN_5399; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_4 <= 1'h0;
      end else begin
        mask_7_2_4 <= _GEN_1351;
      end
    end else begin
      mask_7_2_4 <= _GEN_1351;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_7_2_5 <= _GEN_9559;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_7_2_5 <= _GEN_5463; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_5 <= 1'h0;
      end else begin
        mask_7_2_5 <= _GEN_1367;
      end
    end else begin
      mask_7_2_5 <= _GEN_1367;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_7_2_6 <= _GEN_9623;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_7_2_6 <= _GEN_5527; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_6 <= 1'h0;
      end else begin
        mask_7_2_6 <= _GEN_1383;
      end
    end else begin
      mask_7_2_6 <= _GEN_1383;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_7_2_7 <= _GEN_9687;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_7_2_7 <= _GEN_5591; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_2_7 <= 1'h0;
      end else begin
        mask_7_2_7 <= _GEN_1399;
      end
    end else begin
      mask_7_2_7 <= _GEN_1399;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_7_3_0 <= _GEN_9751;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_7_3_0 <= _GEN_5655; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_0 <= 1'h0;
      end else begin
        mask_7_3_0 <= _GEN_1415;
      end
    end else begin
      mask_7_3_0 <= _GEN_1415;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_7_3_1 <= _GEN_9815;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_7_3_1 <= _GEN_5719; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_1 <= 1'h0;
      end else begin
        mask_7_3_1 <= _GEN_1431;
      end
    end else begin
      mask_7_3_1 <= _GEN_1431;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_7_3_2 <= _GEN_9879;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_7_3_2 <= _GEN_5783; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_2 <= 1'h0;
      end else begin
        mask_7_3_2 <= _GEN_1447;
      end
    end else begin
      mask_7_3_2 <= _GEN_1447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_7_3_3 <= _GEN_9943;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_7_3_3 <= _GEN_5847; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_3 <= 1'h0;
      end else begin
        mask_7_3_3 <= _GEN_1463;
      end
    end else begin
      mask_7_3_3 <= _GEN_1463;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_7_3_4 <= _GEN_10007;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_7_3_4 <= _GEN_5911; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_4 <= 1'h0;
      end else begin
        mask_7_3_4 <= _GEN_1479;
      end
    end else begin
      mask_7_3_4 <= _GEN_1479;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_7_3_5 <= _GEN_10071;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_7_3_5 <= _GEN_5975; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_5 <= 1'h0;
      end else begin
        mask_7_3_5 <= _GEN_1495;
      end
    end else begin
      mask_7_3_5 <= _GEN_1495;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_7_3_6 <= _GEN_10135;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_7_3_6 <= _GEN_6039; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_6 <= 1'h0;
      end else begin
        mask_7_3_6 <= _GEN_1511;
      end
    end else begin
      mask_7_3_6 <= _GEN_1511;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_7_3_7 <= _GEN_10199;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_7_3_7 <= _GEN_6103; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_3_7 <= 1'h0;
      end else begin
        mask_7_3_7 <= _GEN_1527;
      end
    end else begin
      mask_7_3_7 <= _GEN_1527;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_7_4_0 <= _GEN_10263;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_7_4_0 <= _GEN_6167; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_0 <= 1'h0;
      end else begin
        mask_7_4_0 <= _GEN_1543;
      end
    end else begin
      mask_7_4_0 <= _GEN_1543;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_7_4_1 <= _GEN_10327;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_7_4_1 <= _GEN_6231; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_1 <= 1'h0;
      end else begin
        mask_7_4_1 <= _GEN_1559;
      end
    end else begin
      mask_7_4_1 <= _GEN_1559;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_7_4_2 <= _GEN_10391;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_7_4_2 <= _GEN_6295; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_2 <= 1'h0;
      end else begin
        mask_7_4_2 <= _GEN_1575;
      end
    end else begin
      mask_7_4_2 <= _GEN_1575;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_7_4_3 <= _GEN_10455;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_7_4_3 <= _GEN_6359; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_3 <= 1'h0;
      end else begin
        mask_7_4_3 <= _GEN_1591;
      end
    end else begin
      mask_7_4_3 <= _GEN_1591;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_7_4_4 <= _GEN_10519;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_7_4_4 <= _GEN_6423; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_4 <= 1'h0;
      end else begin
        mask_7_4_4 <= _GEN_1607;
      end
    end else begin
      mask_7_4_4 <= _GEN_1607;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_7_4_5 <= _GEN_10583;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_7_4_5 <= _GEN_6487; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_5 <= 1'h0;
      end else begin
        mask_7_4_5 <= _GEN_1623;
      end
    end else begin
      mask_7_4_5 <= _GEN_1623;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_7_4_6 <= _GEN_10647;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_7_4_6 <= _GEN_6551; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_6 <= 1'h0;
      end else begin
        mask_7_4_6 <= _GEN_1639;
      end
    end else begin
      mask_7_4_6 <= _GEN_1639;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_7_4_7 <= _GEN_10711;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_7_4_7 <= _GEN_6615; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_4_7 <= 1'h0;
      end else begin
        mask_7_4_7 <= _GEN_1655;
      end
    end else begin
      mask_7_4_7 <= _GEN_1655;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_7_5_0 <= _GEN_10775;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_7_5_0 <= _GEN_6679; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_0 <= 1'h0;
      end else begin
        mask_7_5_0 <= _GEN_1671;
      end
    end else begin
      mask_7_5_0 <= _GEN_1671;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_7_5_1 <= _GEN_10839;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_7_5_1 <= _GEN_6743; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_1 <= 1'h0;
      end else begin
        mask_7_5_1 <= _GEN_1687;
      end
    end else begin
      mask_7_5_1 <= _GEN_1687;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_7_5_2 <= _GEN_10903;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_7_5_2 <= _GEN_6807; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_2 <= 1'h0;
      end else begin
        mask_7_5_2 <= _GEN_1703;
      end
    end else begin
      mask_7_5_2 <= _GEN_1703;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_7_5_3 <= _GEN_10967;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_7_5_3 <= _GEN_6871; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_3 <= 1'h0;
      end else begin
        mask_7_5_3 <= _GEN_1719;
      end
    end else begin
      mask_7_5_3 <= _GEN_1719;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_7_5_4 <= _GEN_11031;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_7_5_4 <= _GEN_6935; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_4 <= 1'h0;
      end else begin
        mask_7_5_4 <= _GEN_1735;
      end
    end else begin
      mask_7_5_4 <= _GEN_1735;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_7_5_5 <= _GEN_11095;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_7_5_5 <= _GEN_6999; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_5 <= 1'h0;
      end else begin
        mask_7_5_5 <= _GEN_1751;
      end
    end else begin
      mask_7_5_5 <= _GEN_1751;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_7_5_6 <= _GEN_11159;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_7_5_6 <= _GEN_7063; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_6 <= 1'h0;
      end else begin
        mask_7_5_6 <= _GEN_1767;
      end
    end else begin
      mask_7_5_6 <= _GEN_1767;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_7_5_7 <= _GEN_11223;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_7_5_7 <= _GEN_7127; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_5_7 <= 1'h0;
      end else begin
        mask_7_5_7 <= _GEN_1783;
      end
    end else begin
      mask_7_5_7 <= _GEN_1783;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_7_6_0 <= _GEN_11287;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_7_6_0 <= _GEN_7191; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_0 <= 1'h0;
      end else begin
        mask_7_6_0 <= _GEN_1799;
      end
    end else begin
      mask_7_6_0 <= _GEN_1799;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_7_6_1 <= _GEN_11351;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_7_6_1 <= _GEN_7255; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_1 <= 1'h0;
      end else begin
        mask_7_6_1 <= _GEN_1815;
      end
    end else begin
      mask_7_6_1 <= _GEN_1815;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_7_6_2 <= _GEN_11415;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_7_6_2 <= _GEN_7319; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_2 <= 1'h0;
      end else begin
        mask_7_6_2 <= _GEN_1831;
      end
    end else begin
      mask_7_6_2 <= _GEN_1831;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_7_6_3 <= _GEN_11479;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_7_6_3 <= _GEN_7383; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_3 <= 1'h0;
      end else begin
        mask_7_6_3 <= _GEN_1847;
      end
    end else begin
      mask_7_6_3 <= _GEN_1847;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_7_6_4 <= _GEN_11543;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_7_6_4 <= _GEN_7447; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_4 <= 1'h0;
      end else begin
        mask_7_6_4 <= _GEN_1863;
      end
    end else begin
      mask_7_6_4 <= _GEN_1863;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_7_6_5 <= _GEN_11607;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_7_6_5 <= _GEN_7511; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_5 <= 1'h0;
      end else begin
        mask_7_6_5 <= _GEN_1879;
      end
    end else begin
      mask_7_6_5 <= _GEN_1879;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_7_6_6 <= _GEN_11671;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_7_6_6 <= _GEN_7575; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_6 <= 1'h0;
      end else begin
        mask_7_6_6 <= _GEN_1895;
      end
    end else begin
      mask_7_6_6 <= _GEN_1895;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_7_6_7 <= _GEN_11735;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_7_6_7 <= _GEN_7639; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_6_7 <= 1'h0;
      end else begin
        mask_7_6_7 <= _GEN_1911;
      end
    end else begin
      mask_7_6_7 <= _GEN_1911;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_7_7_0 <= _GEN_11799;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_7_7_0 <= _GEN_7703; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_0 <= 1'h0;
      end else begin
        mask_7_7_0 <= _GEN_1927;
      end
    end else begin
      mask_7_7_0 <= _GEN_1927;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_7_7_1 <= _GEN_11863;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_7_7_1 <= _GEN_7767; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_1 <= 1'h0;
      end else begin
        mask_7_7_1 <= _GEN_1943;
      end
    end else begin
      mask_7_7_1 <= _GEN_1943;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_7_7_2 <= _GEN_11927;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_7_7_2 <= _GEN_7831; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_2 <= 1'h0;
      end else begin
        mask_7_7_2 <= _GEN_1959;
      end
    end else begin
      mask_7_7_2 <= _GEN_1959;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_7_7_3 <= _GEN_11991;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_7_7_3 <= _GEN_7895; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_3 <= 1'h0;
      end else begin
        mask_7_7_3 <= _GEN_1975;
      end
    end else begin
      mask_7_7_3 <= _GEN_1975;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_7_7_4 <= _GEN_12055;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_7_7_4 <= _GEN_7959; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_4 <= 1'h0;
      end else begin
        mask_7_7_4 <= _GEN_1991;
      end
    end else begin
      mask_7_7_4 <= _GEN_1991;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_7_7_5 <= _GEN_12119;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_7_7_5 <= _GEN_8023; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_5 <= 1'h0;
      end else begin
        mask_7_7_5 <= _GEN_2007;
      end
    end else begin
      mask_7_7_5 <= _GEN_2007;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_7_7_6 <= _GEN_12183;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_7_7_6 <= _GEN_8087; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_6 <= 1'h0;
      end else begin
        mask_7_7_6 <= _GEN_2023;
      end
    end else begin
      mask_7_7_6 <= _GEN_2023;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_7_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_7_7_7 <= _GEN_12247;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_7_7_7 <= _GEN_8151; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h7 == line_mask_clean_line_1) begin
        mask_7_7_7 <= 1'h0;
      end else begin
        mask_7_7_7 <= _GEN_2039;
      end
    end else begin
      mask_7_7_7 <= _GEN_2039;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_8_0_0 <= _GEN_8216;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_8_0_0 <= _GEN_4120; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_0 <= 1'h0;
      end else begin
        mask_8_0_0 <= _GEN_1032;
      end
    end else begin
      mask_8_0_0 <= _GEN_1032;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_8_0_1 <= _GEN_8280;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_8_0_1 <= _GEN_4184; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_1 <= 1'h0;
      end else begin
        mask_8_0_1 <= _GEN_1048;
      end
    end else begin
      mask_8_0_1 <= _GEN_1048;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_8_0_2 <= _GEN_8344;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_8_0_2 <= _GEN_4248; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_2 <= 1'h0;
      end else begin
        mask_8_0_2 <= _GEN_1064;
      end
    end else begin
      mask_8_0_2 <= _GEN_1064;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_8_0_3 <= _GEN_8408;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_8_0_3 <= _GEN_4312; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_3 <= 1'h0;
      end else begin
        mask_8_0_3 <= _GEN_1080;
      end
    end else begin
      mask_8_0_3 <= _GEN_1080;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_8_0_4 <= _GEN_8472;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_8_0_4 <= _GEN_4376; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_4 <= 1'h0;
      end else begin
        mask_8_0_4 <= _GEN_1096;
      end
    end else begin
      mask_8_0_4 <= _GEN_1096;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_8_0_5 <= _GEN_8536;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_8_0_5 <= _GEN_4440; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_5 <= 1'h0;
      end else begin
        mask_8_0_5 <= _GEN_1112;
      end
    end else begin
      mask_8_0_5 <= _GEN_1112;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_8_0_6 <= _GEN_8600;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_8_0_6 <= _GEN_4504; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_6 <= 1'h0;
      end else begin
        mask_8_0_6 <= _GEN_1128;
      end
    end else begin
      mask_8_0_6 <= _GEN_1128;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_8_0_7 <= _GEN_8664;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_8_0_7 <= _GEN_4568; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_0_7 <= 1'h0;
      end else begin
        mask_8_0_7 <= _GEN_1144;
      end
    end else begin
      mask_8_0_7 <= _GEN_1144;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_8_1_0 <= _GEN_8728;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_8_1_0 <= _GEN_4632; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_0 <= 1'h0;
      end else begin
        mask_8_1_0 <= _GEN_1160;
      end
    end else begin
      mask_8_1_0 <= _GEN_1160;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_8_1_1 <= _GEN_8792;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_8_1_1 <= _GEN_4696; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_1 <= 1'h0;
      end else begin
        mask_8_1_1 <= _GEN_1176;
      end
    end else begin
      mask_8_1_1 <= _GEN_1176;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_8_1_2 <= _GEN_8856;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_8_1_2 <= _GEN_4760; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_2 <= 1'h0;
      end else begin
        mask_8_1_2 <= _GEN_1192;
      end
    end else begin
      mask_8_1_2 <= _GEN_1192;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_8_1_3 <= _GEN_8920;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_8_1_3 <= _GEN_4824; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_3 <= 1'h0;
      end else begin
        mask_8_1_3 <= _GEN_1208;
      end
    end else begin
      mask_8_1_3 <= _GEN_1208;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_8_1_4 <= _GEN_8984;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_8_1_4 <= _GEN_4888; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_4 <= 1'h0;
      end else begin
        mask_8_1_4 <= _GEN_1224;
      end
    end else begin
      mask_8_1_4 <= _GEN_1224;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_8_1_5 <= _GEN_9048;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_8_1_5 <= _GEN_4952; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_5 <= 1'h0;
      end else begin
        mask_8_1_5 <= _GEN_1240;
      end
    end else begin
      mask_8_1_5 <= _GEN_1240;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_8_1_6 <= _GEN_9112;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_8_1_6 <= _GEN_5016; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_6 <= 1'h0;
      end else begin
        mask_8_1_6 <= _GEN_1256;
      end
    end else begin
      mask_8_1_6 <= _GEN_1256;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_8_1_7 <= _GEN_9176;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_8_1_7 <= _GEN_5080; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_1_7 <= 1'h0;
      end else begin
        mask_8_1_7 <= _GEN_1272;
      end
    end else begin
      mask_8_1_7 <= _GEN_1272;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_8_2_0 <= _GEN_9240;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_8_2_0 <= _GEN_5144; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_0 <= 1'h0;
      end else begin
        mask_8_2_0 <= _GEN_1288;
      end
    end else begin
      mask_8_2_0 <= _GEN_1288;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_8_2_1 <= _GEN_9304;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_8_2_1 <= _GEN_5208; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_1 <= 1'h0;
      end else begin
        mask_8_2_1 <= _GEN_1304;
      end
    end else begin
      mask_8_2_1 <= _GEN_1304;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_8_2_2 <= _GEN_9368;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_8_2_2 <= _GEN_5272; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_2 <= 1'h0;
      end else begin
        mask_8_2_2 <= _GEN_1320;
      end
    end else begin
      mask_8_2_2 <= _GEN_1320;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_8_2_3 <= _GEN_9432;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_8_2_3 <= _GEN_5336; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_3 <= 1'h0;
      end else begin
        mask_8_2_3 <= _GEN_1336;
      end
    end else begin
      mask_8_2_3 <= _GEN_1336;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_8_2_4 <= _GEN_9496;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_8_2_4 <= _GEN_5400; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_4 <= 1'h0;
      end else begin
        mask_8_2_4 <= _GEN_1352;
      end
    end else begin
      mask_8_2_4 <= _GEN_1352;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_8_2_5 <= _GEN_9560;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_8_2_5 <= _GEN_5464; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_5 <= 1'h0;
      end else begin
        mask_8_2_5 <= _GEN_1368;
      end
    end else begin
      mask_8_2_5 <= _GEN_1368;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_8_2_6 <= _GEN_9624;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_8_2_6 <= _GEN_5528; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_6 <= 1'h0;
      end else begin
        mask_8_2_6 <= _GEN_1384;
      end
    end else begin
      mask_8_2_6 <= _GEN_1384;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_8_2_7 <= _GEN_9688;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_8_2_7 <= _GEN_5592; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_2_7 <= 1'h0;
      end else begin
        mask_8_2_7 <= _GEN_1400;
      end
    end else begin
      mask_8_2_7 <= _GEN_1400;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_8_3_0 <= _GEN_9752;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_8_3_0 <= _GEN_5656; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_0 <= 1'h0;
      end else begin
        mask_8_3_0 <= _GEN_1416;
      end
    end else begin
      mask_8_3_0 <= _GEN_1416;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_8_3_1 <= _GEN_9816;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_8_3_1 <= _GEN_5720; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_1 <= 1'h0;
      end else begin
        mask_8_3_1 <= _GEN_1432;
      end
    end else begin
      mask_8_3_1 <= _GEN_1432;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_8_3_2 <= _GEN_9880;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_8_3_2 <= _GEN_5784; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_2 <= 1'h0;
      end else begin
        mask_8_3_2 <= _GEN_1448;
      end
    end else begin
      mask_8_3_2 <= _GEN_1448;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_8_3_3 <= _GEN_9944;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_8_3_3 <= _GEN_5848; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_3 <= 1'h0;
      end else begin
        mask_8_3_3 <= _GEN_1464;
      end
    end else begin
      mask_8_3_3 <= _GEN_1464;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_8_3_4 <= _GEN_10008;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_8_3_4 <= _GEN_5912; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_4 <= 1'h0;
      end else begin
        mask_8_3_4 <= _GEN_1480;
      end
    end else begin
      mask_8_3_4 <= _GEN_1480;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_8_3_5 <= _GEN_10072;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_8_3_5 <= _GEN_5976; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_5 <= 1'h0;
      end else begin
        mask_8_3_5 <= _GEN_1496;
      end
    end else begin
      mask_8_3_5 <= _GEN_1496;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_8_3_6 <= _GEN_10136;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_8_3_6 <= _GEN_6040; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_6 <= 1'h0;
      end else begin
        mask_8_3_6 <= _GEN_1512;
      end
    end else begin
      mask_8_3_6 <= _GEN_1512;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_8_3_7 <= _GEN_10200;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_8_3_7 <= _GEN_6104; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_3_7 <= 1'h0;
      end else begin
        mask_8_3_7 <= _GEN_1528;
      end
    end else begin
      mask_8_3_7 <= _GEN_1528;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_8_4_0 <= _GEN_10264;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_8_4_0 <= _GEN_6168; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_0 <= 1'h0;
      end else begin
        mask_8_4_0 <= _GEN_1544;
      end
    end else begin
      mask_8_4_0 <= _GEN_1544;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_8_4_1 <= _GEN_10328;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_8_4_1 <= _GEN_6232; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_1 <= 1'h0;
      end else begin
        mask_8_4_1 <= _GEN_1560;
      end
    end else begin
      mask_8_4_1 <= _GEN_1560;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_8_4_2 <= _GEN_10392;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_8_4_2 <= _GEN_6296; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_2 <= 1'h0;
      end else begin
        mask_8_4_2 <= _GEN_1576;
      end
    end else begin
      mask_8_4_2 <= _GEN_1576;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_8_4_3 <= _GEN_10456;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_8_4_3 <= _GEN_6360; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_3 <= 1'h0;
      end else begin
        mask_8_4_3 <= _GEN_1592;
      end
    end else begin
      mask_8_4_3 <= _GEN_1592;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_8_4_4 <= _GEN_10520;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_8_4_4 <= _GEN_6424; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_4 <= 1'h0;
      end else begin
        mask_8_4_4 <= _GEN_1608;
      end
    end else begin
      mask_8_4_4 <= _GEN_1608;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_8_4_5 <= _GEN_10584;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_8_4_5 <= _GEN_6488; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_5 <= 1'h0;
      end else begin
        mask_8_4_5 <= _GEN_1624;
      end
    end else begin
      mask_8_4_5 <= _GEN_1624;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_8_4_6 <= _GEN_10648;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_8_4_6 <= _GEN_6552; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_6 <= 1'h0;
      end else begin
        mask_8_4_6 <= _GEN_1640;
      end
    end else begin
      mask_8_4_6 <= _GEN_1640;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_8_4_7 <= _GEN_10712;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_8_4_7 <= _GEN_6616; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_4_7 <= 1'h0;
      end else begin
        mask_8_4_7 <= _GEN_1656;
      end
    end else begin
      mask_8_4_7 <= _GEN_1656;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_8_5_0 <= _GEN_10776;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_8_5_0 <= _GEN_6680; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_0 <= 1'h0;
      end else begin
        mask_8_5_0 <= _GEN_1672;
      end
    end else begin
      mask_8_5_0 <= _GEN_1672;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_8_5_1 <= _GEN_10840;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_8_5_1 <= _GEN_6744; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_1 <= 1'h0;
      end else begin
        mask_8_5_1 <= _GEN_1688;
      end
    end else begin
      mask_8_5_1 <= _GEN_1688;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_8_5_2 <= _GEN_10904;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_8_5_2 <= _GEN_6808; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_2 <= 1'h0;
      end else begin
        mask_8_5_2 <= _GEN_1704;
      end
    end else begin
      mask_8_5_2 <= _GEN_1704;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_8_5_3 <= _GEN_10968;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_8_5_3 <= _GEN_6872; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_3 <= 1'h0;
      end else begin
        mask_8_5_3 <= _GEN_1720;
      end
    end else begin
      mask_8_5_3 <= _GEN_1720;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_8_5_4 <= _GEN_11032;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_8_5_4 <= _GEN_6936; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_4 <= 1'h0;
      end else begin
        mask_8_5_4 <= _GEN_1736;
      end
    end else begin
      mask_8_5_4 <= _GEN_1736;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_8_5_5 <= _GEN_11096;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_8_5_5 <= _GEN_7000; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_5 <= 1'h0;
      end else begin
        mask_8_5_5 <= _GEN_1752;
      end
    end else begin
      mask_8_5_5 <= _GEN_1752;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_8_5_6 <= _GEN_11160;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_8_5_6 <= _GEN_7064; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_6 <= 1'h0;
      end else begin
        mask_8_5_6 <= _GEN_1768;
      end
    end else begin
      mask_8_5_6 <= _GEN_1768;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_8_5_7 <= _GEN_11224;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_8_5_7 <= _GEN_7128; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_5_7 <= 1'h0;
      end else begin
        mask_8_5_7 <= _GEN_1784;
      end
    end else begin
      mask_8_5_7 <= _GEN_1784;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_8_6_0 <= _GEN_11288;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_8_6_0 <= _GEN_7192; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_0 <= 1'h0;
      end else begin
        mask_8_6_0 <= _GEN_1800;
      end
    end else begin
      mask_8_6_0 <= _GEN_1800;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_8_6_1 <= _GEN_11352;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_8_6_1 <= _GEN_7256; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_1 <= 1'h0;
      end else begin
        mask_8_6_1 <= _GEN_1816;
      end
    end else begin
      mask_8_6_1 <= _GEN_1816;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_8_6_2 <= _GEN_11416;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_8_6_2 <= _GEN_7320; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_2 <= 1'h0;
      end else begin
        mask_8_6_2 <= _GEN_1832;
      end
    end else begin
      mask_8_6_2 <= _GEN_1832;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_8_6_3 <= _GEN_11480;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_8_6_3 <= _GEN_7384; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_3 <= 1'h0;
      end else begin
        mask_8_6_3 <= _GEN_1848;
      end
    end else begin
      mask_8_6_3 <= _GEN_1848;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_8_6_4 <= _GEN_11544;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_8_6_4 <= _GEN_7448; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_4 <= 1'h0;
      end else begin
        mask_8_6_4 <= _GEN_1864;
      end
    end else begin
      mask_8_6_4 <= _GEN_1864;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_8_6_5 <= _GEN_11608;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_8_6_5 <= _GEN_7512; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_5 <= 1'h0;
      end else begin
        mask_8_6_5 <= _GEN_1880;
      end
    end else begin
      mask_8_6_5 <= _GEN_1880;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_8_6_6 <= _GEN_11672;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_8_6_6 <= _GEN_7576; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_6 <= 1'h0;
      end else begin
        mask_8_6_6 <= _GEN_1896;
      end
    end else begin
      mask_8_6_6 <= _GEN_1896;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_8_6_7 <= _GEN_11736;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_8_6_7 <= _GEN_7640; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_6_7 <= 1'h0;
      end else begin
        mask_8_6_7 <= _GEN_1912;
      end
    end else begin
      mask_8_6_7 <= _GEN_1912;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_8_7_0 <= _GEN_11800;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_8_7_0 <= _GEN_7704; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_0 <= 1'h0;
      end else begin
        mask_8_7_0 <= _GEN_1928;
      end
    end else begin
      mask_8_7_0 <= _GEN_1928;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_8_7_1 <= _GEN_11864;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_8_7_1 <= _GEN_7768; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_1 <= 1'h0;
      end else begin
        mask_8_7_1 <= _GEN_1944;
      end
    end else begin
      mask_8_7_1 <= _GEN_1944;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_8_7_2 <= _GEN_11928;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_8_7_2 <= _GEN_7832; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_2 <= 1'h0;
      end else begin
        mask_8_7_2 <= _GEN_1960;
      end
    end else begin
      mask_8_7_2 <= _GEN_1960;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_8_7_3 <= _GEN_11992;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_8_7_3 <= _GEN_7896; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_3 <= 1'h0;
      end else begin
        mask_8_7_3 <= _GEN_1976;
      end
    end else begin
      mask_8_7_3 <= _GEN_1976;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_8_7_4 <= _GEN_12056;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_8_7_4 <= _GEN_7960; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_4 <= 1'h0;
      end else begin
        mask_8_7_4 <= _GEN_1992;
      end
    end else begin
      mask_8_7_4 <= _GEN_1992;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_8_7_5 <= _GEN_12120;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_8_7_5 <= _GEN_8024; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_5 <= 1'h0;
      end else begin
        mask_8_7_5 <= _GEN_2008;
      end
    end else begin
      mask_8_7_5 <= _GEN_2008;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_8_7_6 <= _GEN_12184;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_8_7_6 <= _GEN_8088; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_6 <= 1'h0;
      end else begin
        mask_8_7_6 <= _GEN_2024;
      end
    end else begin
      mask_8_7_6 <= _GEN_2024;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_8_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_8_7_7 <= _GEN_12248;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_8_7_7 <= _GEN_8152; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h8 == line_mask_clean_line_1) begin
        mask_8_7_7 <= 1'h0;
      end else begin
        mask_8_7_7 <= _GEN_2040;
      end
    end else begin
      mask_8_7_7 <= _GEN_2040;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_9_0_0 <= _GEN_8217;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_9_0_0 <= _GEN_4121; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_0 <= 1'h0;
      end else begin
        mask_9_0_0 <= _GEN_1033;
      end
    end else begin
      mask_9_0_0 <= _GEN_1033;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_9_0_1 <= _GEN_8281;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_9_0_1 <= _GEN_4185; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_1 <= 1'h0;
      end else begin
        mask_9_0_1 <= _GEN_1049;
      end
    end else begin
      mask_9_0_1 <= _GEN_1049;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_9_0_2 <= _GEN_8345;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_9_0_2 <= _GEN_4249; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_2 <= 1'h0;
      end else begin
        mask_9_0_2 <= _GEN_1065;
      end
    end else begin
      mask_9_0_2 <= _GEN_1065;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_9_0_3 <= _GEN_8409;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_9_0_3 <= _GEN_4313; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_3 <= 1'h0;
      end else begin
        mask_9_0_3 <= _GEN_1081;
      end
    end else begin
      mask_9_0_3 <= _GEN_1081;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_9_0_4 <= _GEN_8473;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_9_0_4 <= _GEN_4377; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_4 <= 1'h0;
      end else begin
        mask_9_0_4 <= _GEN_1097;
      end
    end else begin
      mask_9_0_4 <= _GEN_1097;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_9_0_5 <= _GEN_8537;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_9_0_5 <= _GEN_4441; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_5 <= 1'h0;
      end else begin
        mask_9_0_5 <= _GEN_1113;
      end
    end else begin
      mask_9_0_5 <= _GEN_1113;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_9_0_6 <= _GEN_8601;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_9_0_6 <= _GEN_4505; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_6 <= 1'h0;
      end else begin
        mask_9_0_6 <= _GEN_1129;
      end
    end else begin
      mask_9_0_6 <= _GEN_1129;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_9_0_7 <= _GEN_8665;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_9_0_7 <= _GEN_4569; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_0_7 <= 1'h0;
      end else begin
        mask_9_0_7 <= _GEN_1145;
      end
    end else begin
      mask_9_0_7 <= _GEN_1145;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_9_1_0 <= _GEN_8729;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_9_1_0 <= _GEN_4633; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_0 <= 1'h0;
      end else begin
        mask_9_1_0 <= _GEN_1161;
      end
    end else begin
      mask_9_1_0 <= _GEN_1161;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_9_1_1 <= _GEN_8793;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_9_1_1 <= _GEN_4697; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_1 <= 1'h0;
      end else begin
        mask_9_1_1 <= _GEN_1177;
      end
    end else begin
      mask_9_1_1 <= _GEN_1177;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_9_1_2 <= _GEN_8857;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_9_1_2 <= _GEN_4761; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_2 <= 1'h0;
      end else begin
        mask_9_1_2 <= _GEN_1193;
      end
    end else begin
      mask_9_1_2 <= _GEN_1193;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_9_1_3 <= _GEN_8921;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_9_1_3 <= _GEN_4825; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_3 <= 1'h0;
      end else begin
        mask_9_1_3 <= _GEN_1209;
      end
    end else begin
      mask_9_1_3 <= _GEN_1209;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_9_1_4 <= _GEN_8985;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_9_1_4 <= _GEN_4889; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_4 <= 1'h0;
      end else begin
        mask_9_1_4 <= _GEN_1225;
      end
    end else begin
      mask_9_1_4 <= _GEN_1225;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_9_1_5 <= _GEN_9049;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_9_1_5 <= _GEN_4953; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_5 <= 1'h0;
      end else begin
        mask_9_1_5 <= _GEN_1241;
      end
    end else begin
      mask_9_1_5 <= _GEN_1241;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_9_1_6 <= _GEN_9113;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_9_1_6 <= _GEN_5017; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_6 <= 1'h0;
      end else begin
        mask_9_1_6 <= _GEN_1257;
      end
    end else begin
      mask_9_1_6 <= _GEN_1257;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_9_1_7 <= _GEN_9177;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_9_1_7 <= _GEN_5081; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_1_7 <= 1'h0;
      end else begin
        mask_9_1_7 <= _GEN_1273;
      end
    end else begin
      mask_9_1_7 <= _GEN_1273;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_9_2_0 <= _GEN_9241;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_9_2_0 <= _GEN_5145; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_0 <= 1'h0;
      end else begin
        mask_9_2_0 <= _GEN_1289;
      end
    end else begin
      mask_9_2_0 <= _GEN_1289;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_9_2_1 <= _GEN_9305;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_9_2_1 <= _GEN_5209; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_1 <= 1'h0;
      end else begin
        mask_9_2_1 <= _GEN_1305;
      end
    end else begin
      mask_9_2_1 <= _GEN_1305;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_9_2_2 <= _GEN_9369;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_9_2_2 <= _GEN_5273; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_2 <= 1'h0;
      end else begin
        mask_9_2_2 <= _GEN_1321;
      end
    end else begin
      mask_9_2_2 <= _GEN_1321;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_9_2_3 <= _GEN_9433;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_9_2_3 <= _GEN_5337; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_3 <= 1'h0;
      end else begin
        mask_9_2_3 <= _GEN_1337;
      end
    end else begin
      mask_9_2_3 <= _GEN_1337;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_9_2_4 <= _GEN_9497;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_9_2_4 <= _GEN_5401; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_4 <= 1'h0;
      end else begin
        mask_9_2_4 <= _GEN_1353;
      end
    end else begin
      mask_9_2_4 <= _GEN_1353;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_9_2_5 <= _GEN_9561;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_9_2_5 <= _GEN_5465; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_5 <= 1'h0;
      end else begin
        mask_9_2_5 <= _GEN_1369;
      end
    end else begin
      mask_9_2_5 <= _GEN_1369;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_9_2_6 <= _GEN_9625;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_9_2_6 <= _GEN_5529; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_6 <= 1'h0;
      end else begin
        mask_9_2_6 <= _GEN_1385;
      end
    end else begin
      mask_9_2_6 <= _GEN_1385;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_9_2_7 <= _GEN_9689;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_9_2_7 <= _GEN_5593; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_2_7 <= 1'h0;
      end else begin
        mask_9_2_7 <= _GEN_1401;
      end
    end else begin
      mask_9_2_7 <= _GEN_1401;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_9_3_0 <= _GEN_9753;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_9_3_0 <= _GEN_5657; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_0 <= 1'h0;
      end else begin
        mask_9_3_0 <= _GEN_1417;
      end
    end else begin
      mask_9_3_0 <= _GEN_1417;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_9_3_1 <= _GEN_9817;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_9_3_1 <= _GEN_5721; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_1 <= 1'h0;
      end else begin
        mask_9_3_1 <= _GEN_1433;
      end
    end else begin
      mask_9_3_1 <= _GEN_1433;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_9_3_2 <= _GEN_9881;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_9_3_2 <= _GEN_5785; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_2 <= 1'h0;
      end else begin
        mask_9_3_2 <= _GEN_1449;
      end
    end else begin
      mask_9_3_2 <= _GEN_1449;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_9_3_3 <= _GEN_9945;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_9_3_3 <= _GEN_5849; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_3 <= 1'h0;
      end else begin
        mask_9_3_3 <= _GEN_1465;
      end
    end else begin
      mask_9_3_3 <= _GEN_1465;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_9_3_4 <= _GEN_10009;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_9_3_4 <= _GEN_5913; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_4 <= 1'h0;
      end else begin
        mask_9_3_4 <= _GEN_1481;
      end
    end else begin
      mask_9_3_4 <= _GEN_1481;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_9_3_5 <= _GEN_10073;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_9_3_5 <= _GEN_5977; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_5 <= 1'h0;
      end else begin
        mask_9_3_5 <= _GEN_1497;
      end
    end else begin
      mask_9_3_5 <= _GEN_1497;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_9_3_6 <= _GEN_10137;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_9_3_6 <= _GEN_6041; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_6 <= 1'h0;
      end else begin
        mask_9_3_6 <= _GEN_1513;
      end
    end else begin
      mask_9_3_6 <= _GEN_1513;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_9_3_7 <= _GEN_10201;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_9_3_7 <= _GEN_6105; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_3_7 <= 1'h0;
      end else begin
        mask_9_3_7 <= _GEN_1529;
      end
    end else begin
      mask_9_3_7 <= _GEN_1529;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_9_4_0 <= _GEN_10265;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_9_4_0 <= _GEN_6169; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_0 <= 1'h0;
      end else begin
        mask_9_4_0 <= _GEN_1545;
      end
    end else begin
      mask_9_4_0 <= _GEN_1545;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_9_4_1 <= _GEN_10329;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_9_4_1 <= _GEN_6233; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_1 <= 1'h0;
      end else begin
        mask_9_4_1 <= _GEN_1561;
      end
    end else begin
      mask_9_4_1 <= _GEN_1561;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_9_4_2 <= _GEN_10393;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_9_4_2 <= _GEN_6297; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_2 <= 1'h0;
      end else begin
        mask_9_4_2 <= _GEN_1577;
      end
    end else begin
      mask_9_4_2 <= _GEN_1577;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_9_4_3 <= _GEN_10457;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_9_4_3 <= _GEN_6361; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_3 <= 1'h0;
      end else begin
        mask_9_4_3 <= _GEN_1593;
      end
    end else begin
      mask_9_4_3 <= _GEN_1593;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_9_4_4 <= _GEN_10521;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_9_4_4 <= _GEN_6425; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_4 <= 1'h0;
      end else begin
        mask_9_4_4 <= _GEN_1609;
      end
    end else begin
      mask_9_4_4 <= _GEN_1609;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_9_4_5 <= _GEN_10585;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_9_4_5 <= _GEN_6489; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_5 <= 1'h0;
      end else begin
        mask_9_4_5 <= _GEN_1625;
      end
    end else begin
      mask_9_4_5 <= _GEN_1625;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_9_4_6 <= _GEN_10649;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_9_4_6 <= _GEN_6553; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_6 <= 1'h0;
      end else begin
        mask_9_4_6 <= _GEN_1641;
      end
    end else begin
      mask_9_4_6 <= _GEN_1641;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_9_4_7 <= _GEN_10713;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_9_4_7 <= _GEN_6617; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_4_7 <= 1'h0;
      end else begin
        mask_9_4_7 <= _GEN_1657;
      end
    end else begin
      mask_9_4_7 <= _GEN_1657;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_9_5_0 <= _GEN_10777;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_9_5_0 <= _GEN_6681; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_0 <= 1'h0;
      end else begin
        mask_9_5_0 <= _GEN_1673;
      end
    end else begin
      mask_9_5_0 <= _GEN_1673;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_9_5_1 <= _GEN_10841;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_9_5_1 <= _GEN_6745; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_1 <= 1'h0;
      end else begin
        mask_9_5_1 <= _GEN_1689;
      end
    end else begin
      mask_9_5_1 <= _GEN_1689;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_9_5_2 <= _GEN_10905;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_9_5_2 <= _GEN_6809; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_2 <= 1'h0;
      end else begin
        mask_9_5_2 <= _GEN_1705;
      end
    end else begin
      mask_9_5_2 <= _GEN_1705;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_9_5_3 <= _GEN_10969;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_9_5_3 <= _GEN_6873; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_3 <= 1'h0;
      end else begin
        mask_9_5_3 <= _GEN_1721;
      end
    end else begin
      mask_9_5_3 <= _GEN_1721;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_9_5_4 <= _GEN_11033;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_9_5_4 <= _GEN_6937; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_4 <= 1'h0;
      end else begin
        mask_9_5_4 <= _GEN_1737;
      end
    end else begin
      mask_9_5_4 <= _GEN_1737;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_9_5_5 <= _GEN_11097;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_9_5_5 <= _GEN_7001; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_5 <= 1'h0;
      end else begin
        mask_9_5_5 <= _GEN_1753;
      end
    end else begin
      mask_9_5_5 <= _GEN_1753;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_9_5_6 <= _GEN_11161;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_9_5_6 <= _GEN_7065; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_6 <= 1'h0;
      end else begin
        mask_9_5_6 <= _GEN_1769;
      end
    end else begin
      mask_9_5_6 <= _GEN_1769;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_9_5_7 <= _GEN_11225;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_9_5_7 <= _GEN_7129; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_5_7 <= 1'h0;
      end else begin
        mask_9_5_7 <= _GEN_1785;
      end
    end else begin
      mask_9_5_7 <= _GEN_1785;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_9_6_0 <= _GEN_11289;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_9_6_0 <= _GEN_7193; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_0 <= 1'h0;
      end else begin
        mask_9_6_0 <= _GEN_1801;
      end
    end else begin
      mask_9_6_0 <= _GEN_1801;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_9_6_1 <= _GEN_11353;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_9_6_1 <= _GEN_7257; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_1 <= 1'h0;
      end else begin
        mask_9_6_1 <= _GEN_1817;
      end
    end else begin
      mask_9_6_1 <= _GEN_1817;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_9_6_2 <= _GEN_11417;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_9_6_2 <= _GEN_7321; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_2 <= 1'h0;
      end else begin
        mask_9_6_2 <= _GEN_1833;
      end
    end else begin
      mask_9_6_2 <= _GEN_1833;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_9_6_3 <= _GEN_11481;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_9_6_3 <= _GEN_7385; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_3 <= 1'h0;
      end else begin
        mask_9_6_3 <= _GEN_1849;
      end
    end else begin
      mask_9_6_3 <= _GEN_1849;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_9_6_4 <= _GEN_11545;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_9_6_4 <= _GEN_7449; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_4 <= 1'h0;
      end else begin
        mask_9_6_4 <= _GEN_1865;
      end
    end else begin
      mask_9_6_4 <= _GEN_1865;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_9_6_5 <= _GEN_11609;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_9_6_5 <= _GEN_7513; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_5 <= 1'h0;
      end else begin
        mask_9_6_5 <= _GEN_1881;
      end
    end else begin
      mask_9_6_5 <= _GEN_1881;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_9_6_6 <= _GEN_11673;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_9_6_6 <= _GEN_7577; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_6 <= 1'h0;
      end else begin
        mask_9_6_6 <= _GEN_1897;
      end
    end else begin
      mask_9_6_6 <= _GEN_1897;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_9_6_7 <= _GEN_11737;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_9_6_7 <= _GEN_7641; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_6_7 <= 1'h0;
      end else begin
        mask_9_6_7 <= _GEN_1913;
      end
    end else begin
      mask_9_6_7 <= _GEN_1913;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_9_7_0 <= _GEN_11801;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_9_7_0 <= _GEN_7705; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_0 <= 1'h0;
      end else begin
        mask_9_7_0 <= _GEN_1929;
      end
    end else begin
      mask_9_7_0 <= _GEN_1929;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_9_7_1 <= _GEN_11865;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_9_7_1 <= _GEN_7769; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_1 <= 1'h0;
      end else begin
        mask_9_7_1 <= _GEN_1945;
      end
    end else begin
      mask_9_7_1 <= _GEN_1945;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_9_7_2 <= _GEN_11929;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_9_7_2 <= _GEN_7833; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_2 <= 1'h0;
      end else begin
        mask_9_7_2 <= _GEN_1961;
      end
    end else begin
      mask_9_7_2 <= _GEN_1961;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_9_7_3 <= _GEN_11993;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_9_7_3 <= _GEN_7897; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_3 <= 1'h0;
      end else begin
        mask_9_7_3 <= _GEN_1977;
      end
    end else begin
      mask_9_7_3 <= _GEN_1977;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_9_7_4 <= _GEN_12057;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_9_7_4 <= _GEN_7961; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_4 <= 1'h0;
      end else begin
        mask_9_7_4 <= _GEN_1993;
      end
    end else begin
      mask_9_7_4 <= _GEN_1993;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_9_7_5 <= _GEN_12121;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_9_7_5 <= _GEN_8025; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_5 <= 1'h0;
      end else begin
        mask_9_7_5 <= _GEN_2009;
      end
    end else begin
      mask_9_7_5 <= _GEN_2009;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_9_7_6 <= _GEN_12185;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_9_7_6 <= _GEN_8089; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_6 <= 1'h0;
      end else begin
        mask_9_7_6 <= _GEN_2025;
      end
    end else begin
      mask_9_7_6 <= _GEN_2025;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_9_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_9_7_7 <= _GEN_12249;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_9_7_7 <= _GEN_8153; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'h9 == line_mask_clean_line_1) begin
        mask_9_7_7 <= 1'h0;
      end else begin
        mask_9_7_7 <= _GEN_2041;
      end
    end else begin
      mask_9_7_7 <= _GEN_2041;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_10_0_0 <= _GEN_8218;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_10_0_0 <= _GEN_4122; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_0 <= 1'h0;
      end else begin
        mask_10_0_0 <= _GEN_1034;
      end
    end else begin
      mask_10_0_0 <= _GEN_1034;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_10_0_1 <= _GEN_8282;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_10_0_1 <= _GEN_4186; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_1 <= 1'h0;
      end else begin
        mask_10_0_1 <= _GEN_1050;
      end
    end else begin
      mask_10_0_1 <= _GEN_1050;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_10_0_2 <= _GEN_8346;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_10_0_2 <= _GEN_4250; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_2 <= 1'h0;
      end else begin
        mask_10_0_2 <= _GEN_1066;
      end
    end else begin
      mask_10_0_2 <= _GEN_1066;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_10_0_3 <= _GEN_8410;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_10_0_3 <= _GEN_4314; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_3 <= 1'h0;
      end else begin
        mask_10_0_3 <= _GEN_1082;
      end
    end else begin
      mask_10_0_3 <= _GEN_1082;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_10_0_4 <= _GEN_8474;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_10_0_4 <= _GEN_4378; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_4 <= 1'h0;
      end else begin
        mask_10_0_4 <= _GEN_1098;
      end
    end else begin
      mask_10_0_4 <= _GEN_1098;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_10_0_5 <= _GEN_8538;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_10_0_5 <= _GEN_4442; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_5 <= 1'h0;
      end else begin
        mask_10_0_5 <= _GEN_1114;
      end
    end else begin
      mask_10_0_5 <= _GEN_1114;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_10_0_6 <= _GEN_8602;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_10_0_6 <= _GEN_4506; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_6 <= 1'h0;
      end else begin
        mask_10_0_6 <= _GEN_1130;
      end
    end else begin
      mask_10_0_6 <= _GEN_1130;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_10_0_7 <= _GEN_8666;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_10_0_7 <= _GEN_4570; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_0_7 <= 1'h0;
      end else begin
        mask_10_0_7 <= _GEN_1146;
      end
    end else begin
      mask_10_0_7 <= _GEN_1146;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_10_1_0 <= _GEN_8730;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_10_1_0 <= _GEN_4634; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_0 <= 1'h0;
      end else begin
        mask_10_1_0 <= _GEN_1162;
      end
    end else begin
      mask_10_1_0 <= _GEN_1162;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_10_1_1 <= _GEN_8794;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_10_1_1 <= _GEN_4698; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_1 <= 1'h0;
      end else begin
        mask_10_1_1 <= _GEN_1178;
      end
    end else begin
      mask_10_1_1 <= _GEN_1178;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_10_1_2 <= _GEN_8858;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_10_1_2 <= _GEN_4762; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_2 <= 1'h0;
      end else begin
        mask_10_1_2 <= _GEN_1194;
      end
    end else begin
      mask_10_1_2 <= _GEN_1194;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_10_1_3 <= _GEN_8922;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_10_1_3 <= _GEN_4826; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_3 <= 1'h0;
      end else begin
        mask_10_1_3 <= _GEN_1210;
      end
    end else begin
      mask_10_1_3 <= _GEN_1210;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_10_1_4 <= _GEN_8986;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_10_1_4 <= _GEN_4890; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_4 <= 1'h0;
      end else begin
        mask_10_1_4 <= _GEN_1226;
      end
    end else begin
      mask_10_1_4 <= _GEN_1226;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_10_1_5 <= _GEN_9050;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_10_1_5 <= _GEN_4954; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_5 <= 1'h0;
      end else begin
        mask_10_1_5 <= _GEN_1242;
      end
    end else begin
      mask_10_1_5 <= _GEN_1242;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_10_1_6 <= _GEN_9114;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_10_1_6 <= _GEN_5018; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_6 <= 1'h0;
      end else begin
        mask_10_1_6 <= _GEN_1258;
      end
    end else begin
      mask_10_1_6 <= _GEN_1258;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_10_1_7 <= _GEN_9178;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_10_1_7 <= _GEN_5082; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_1_7 <= 1'h0;
      end else begin
        mask_10_1_7 <= _GEN_1274;
      end
    end else begin
      mask_10_1_7 <= _GEN_1274;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_10_2_0 <= _GEN_9242;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_10_2_0 <= _GEN_5146; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_0 <= 1'h0;
      end else begin
        mask_10_2_0 <= _GEN_1290;
      end
    end else begin
      mask_10_2_0 <= _GEN_1290;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_10_2_1 <= _GEN_9306;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_10_2_1 <= _GEN_5210; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_1 <= 1'h0;
      end else begin
        mask_10_2_1 <= _GEN_1306;
      end
    end else begin
      mask_10_2_1 <= _GEN_1306;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_10_2_2 <= _GEN_9370;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_10_2_2 <= _GEN_5274; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_2 <= 1'h0;
      end else begin
        mask_10_2_2 <= _GEN_1322;
      end
    end else begin
      mask_10_2_2 <= _GEN_1322;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_10_2_3 <= _GEN_9434;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_10_2_3 <= _GEN_5338; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_3 <= 1'h0;
      end else begin
        mask_10_2_3 <= _GEN_1338;
      end
    end else begin
      mask_10_2_3 <= _GEN_1338;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_10_2_4 <= _GEN_9498;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_10_2_4 <= _GEN_5402; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_4 <= 1'h0;
      end else begin
        mask_10_2_4 <= _GEN_1354;
      end
    end else begin
      mask_10_2_4 <= _GEN_1354;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_10_2_5 <= _GEN_9562;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_10_2_5 <= _GEN_5466; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_5 <= 1'h0;
      end else begin
        mask_10_2_5 <= _GEN_1370;
      end
    end else begin
      mask_10_2_5 <= _GEN_1370;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_10_2_6 <= _GEN_9626;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_10_2_6 <= _GEN_5530; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_6 <= 1'h0;
      end else begin
        mask_10_2_6 <= _GEN_1386;
      end
    end else begin
      mask_10_2_6 <= _GEN_1386;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_10_2_7 <= _GEN_9690;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_10_2_7 <= _GEN_5594; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_2_7 <= 1'h0;
      end else begin
        mask_10_2_7 <= _GEN_1402;
      end
    end else begin
      mask_10_2_7 <= _GEN_1402;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_10_3_0 <= _GEN_9754;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_10_3_0 <= _GEN_5658; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_0 <= 1'h0;
      end else begin
        mask_10_3_0 <= _GEN_1418;
      end
    end else begin
      mask_10_3_0 <= _GEN_1418;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_10_3_1 <= _GEN_9818;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_10_3_1 <= _GEN_5722; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_1 <= 1'h0;
      end else begin
        mask_10_3_1 <= _GEN_1434;
      end
    end else begin
      mask_10_3_1 <= _GEN_1434;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_10_3_2 <= _GEN_9882;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_10_3_2 <= _GEN_5786; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_2 <= 1'h0;
      end else begin
        mask_10_3_2 <= _GEN_1450;
      end
    end else begin
      mask_10_3_2 <= _GEN_1450;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_10_3_3 <= _GEN_9946;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_10_3_3 <= _GEN_5850; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_3 <= 1'h0;
      end else begin
        mask_10_3_3 <= _GEN_1466;
      end
    end else begin
      mask_10_3_3 <= _GEN_1466;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_10_3_4 <= _GEN_10010;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_10_3_4 <= _GEN_5914; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_4 <= 1'h0;
      end else begin
        mask_10_3_4 <= _GEN_1482;
      end
    end else begin
      mask_10_3_4 <= _GEN_1482;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_10_3_5 <= _GEN_10074;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_10_3_5 <= _GEN_5978; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_5 <= 1'h0;
      end else begin
        mask_10_3_5 <= _GEN_1498;
      end
    end else begin
      mask_10_3_5 <= _GEN_1498;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_10_3_6 <= _GEN_10138;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_10_3_6 <= _GEN_6042; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_6 <= 1'h0;
      end else begin
        mask_10_3_6 <= _GEN_1514;
      end
    end else begin
      mask_10_3_6 <= _GEN_1514;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_10_3_7 <= _GEN_10202;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_10_3_7 <= _GEN_6106; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_3_7 <= 1'h0;
      end else begin
        mask_10_3_7 <= _GEN_1530;
      end
    end else begin
      mask_10_3_7 <= _GEN_1530;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_10_4_0 <= _GEN_10266;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_10_4_0 <= _GEN_6170; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_0 <= 1'h0;
      end else begin
        mask_10_4_0 <= _GEN_1546;
      end
    end else begin
      mask_10_4_0 <= _GEN_1546;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_10_4_1 <= _GEN_10330;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_10_4_1 <= _GEN_6234; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_1 <= 1'h0;
      end else begin
        mask_10_4_1 <= _GEN_1562;
      end
    end else begin
      mask_10_4_1 <= _GEN_1562;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_10_4_2 <= _GEN_10394;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_10_4_2 <= _GEN_6298; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_2 <= 1'h0;
      end else begin
        mask_10_4_2 <= _GEN_1578;
      end
    end else begin
      mask_10_4_2 <= _GEN_1578;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_10_4_3 <= _GEN_10458;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_10_4_3 <= _GEN_6362; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_3 <= 1'h0;
      end else begin
        mask_10_4_3 <= _GEN_1594;
      end
    end else begin
      mask_10_4_3 <= _GEN_1594;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_10_4_4 <= _GEN_10522;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_10_4_4 <= _GEN_6426; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_4 <= 1'h0;
      end else begin
        mask_10_4_4 <= _GEN_1610;
      end
    end else begin
      mask_10_4_4 <= _GEN_1610;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_10_4_5 <= _GEN_10586;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_10_4_5 <= _GEN_6490; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_5 <= 1'h0;
      end else begin
        mask_10_4_5 <= _GEN_1626;
      end
    end else begin
      mask_10_4_5 <= _GEN_1626;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_10_4_6 <= _GEN_10650;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_10_4_6 <= _GEN_6554; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_6 <= 1'h0;
      end else begin
        mask_10_4_6 <= _GEN_1642;
      end
    end else begin
      mask_10_4_6 <= _GEN_1642;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_10_4_7 <= _GEN_10714;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_10_4_7 <= _GEN_6618; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_4_7 <= 1'h0;
      end else begin
        mask_10_4_7 <= _GEN_1658;
      end
    end else begin
      mask_10_4_7 <= _GEN_1658;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_10_5_0 <= _GEN_10778;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_10_5_0 <= _GEN_6682; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_0 <= 1'h0;
      end else begin
        mask_10_5_0 <= _GEN_1674;
      end
    end else begin
      mask_10_5_0 <= _GEN_1674;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_10_5_1 <= _GEN_10842;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_10_5_1 <= _GEN_6746; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_1 <= 1'h0;
      end else begin
        mask_10_5_1 <= _GEN_1690;
      end
    end else begin
      mask_10_5_1 <= _GEN_1690;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_10_5_2 <= _GEN_10906;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_10_5_2 <= _GEN_6810; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_2 <= 1'h0;
      end else begin
        mask_10_5_2 <= _GEN_1706;
      end
    end else begin
      mask_10_5_2 <= _GEN_1706;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_10_5_3 <= _GEN_10970;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_10_5_3 <= _GEN_6874; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_3 <= 1'h0;
      end else begin
        mask_10_5_3 <= _GEN_1722;
      end
    end else begin
      mask_10_5_3 <= _GEN_1722;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_10_5_4 <= _GEN_11034;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_10_5_4 <= _GEN_6938; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_4 <= 1'h0;
      end else begin
        mask_10_5_4 <= _GEN_1738;
      end
    end else begin
      mask_10_5_4 <= _GEN_1738;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_10_5_5 <= _GEN_11098;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_10_5_5 <= _GEN_7002; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_5 <= 1'h0;
      end else begin
        mask_10_5_5 <= _GEN_1754;
      end
    end else begin
      mask_10_5_5 <= _GEN_1754;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_10_5_6 <= _GEN_11162;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_10_5_6 <= _GEN_7066; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_6 <= 1'h0;
      end else begin
        mask_10_5_6 <= _GEN_1770;
      end
    end else begin
      mask_10_5_6 <= _GEN_1770;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_10_5_7 <= _GEN_11226;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_10_5_7 <= _GEN_7130; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_5_7 <= 1'h0;
      end else begin
        mask_10_5_7 <= _GEN_1786;
      end
    end else begin
      mask_10_5_7 <= _GEN_1786;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_10_6_0 <= _GEN_11290;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_10_6_0 <= _GEN_7194; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_0 <= 1'h0;
      end else begin
        mask_10_6_0 <= _GEN_1802;
      end
    end else begin
      mask_10_6_0 <= _GEN_1802;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_10_6_1 <= _GEN_11354;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_10_6_1 <= _GEN_7258; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_1 <= 1'h0;
      end else begin
        mask_10_6_1 <= _GEN_1818;
      end
    end else begin
      mask_10_6_1 <= _GEN_1818;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_10_6_2 <= _GEN_11418;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_10_6_2 <= _GEN_7322; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_2 <= 1'h0;
      end else begin
        mask_10_6_2 <= _GEN_1834;
      end
    end else begin
      mask_10_6_2 <= _GEN_1834;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_10_6_3 <= _GEN_11482;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_10_6_3 <= _GEN_7386; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_3 <= 1'h0;
      end else begin
        mask_10_6_3 <= _GEN_1850;
      end
    end else begin
      mask_10_6_3 <= _GEN_1850;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_10_6_4 <= _GEN_11546;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_10_6_4 <= _GEN_7450; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_4 <= 1'h0;
      end else begin
        mask_10_6_4 <= _GEN_1866;
      end
    end else begin
      mask_10_6_4 <= _GEN_1866;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_10_6_5 <= _GEN_11610;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_10_6_5 <= _GEN_7514; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_5 <= 1'h0;
      end else begin
        mask_10_6_5 <= _GEN_1882;
      end
    end else begin
      mask_10_6_5 <= _GEN_1882;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_10_6_6 <= _GEN_11674;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_10_6_6 <= _GEN_7578; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_6 <= 1'h0;
      end else begin
        mask_10_6_6 <= _GEN_1898;
      end
    end else begin
      mask_10_6_6 <= _GEN_1898;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_10_6_7 <= _GEN_11738;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_10_6_7 <= _GEN_7642; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_6_7 <= 1'h0;
      end else begin
        mask_10_6_7 <= _GEN_1914;
      end
    end else begin
      mask_10_6_7 <= _GEN_1914;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_10_7_0 <= _GEN_11802;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_10_7_0 <= _GEN_7706; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_0 <= 1'h0;
      end else begin
        mask_10_7_0 <= _GEN_1930;
      end
    end else begin
      mask_10_7_0 <= _GEN_1930;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_10_7_1 <= _GEN_11866;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_10_7_1 <= _GEN_7770; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_1 <= 1'h0;
      end else begin
        mask_10_7_1 <= _GEN_1946;
      end
    end else begin
      mask_10_7_1 <= _GEN_1946;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_10_7_2 <= _GEN_11930;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_10_7_2 <= _GEN_7834; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_2 <= 1'h0;
      end else begin
        mask_10_7_2 <= _GEN_1962;
      end
    end else begin
      mask_10_7_2 <= _GEN_1962;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_10_7_3 <= _GEN_11994;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_10_7_3 <= _GEN_7898; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_3 <= 1'h0;
      end else begin
        mask_10_7_3 <= _GEN_1978;
      end
    end else begin
      mask_10_7_3 <= _GEN_1978;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_10_7_4 <= _GEN_12058;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_10_7_4 <= _GEN_7962; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_4 <= 1'h0;
      end else begin
        mask_10_7_4 <= _GEN_1994;
      end
    end else begin
      mask_10_7_4 <= _GEN_1994;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_10_7_5 <= _GEN_12122;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_10_7_5 <= _GEN_8026; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_5 <= 1'h0;
      end else begin
        mask_10_7_5 <= _GEN_2010;
      end
    end else begin
      mask_10_7_5 <= _GEN_2010;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_10_7_6 <= _GEN_12186;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_10_7_6 <= _GEN_8090; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_6 <= 1'h0;
      end else begin
        mask_10_7_6 <= _GEN_2026;
      end
    end else begin
      mask_10_7_6 <= _GEN_2026;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_10_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_10_7_7 <= _GEN_12250;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_10_7_7 <= _GEN_8154; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'ha == line_mask_clean_line_1) begin
        mask_10_7_7 <= 1'h0;
      end else begin
        mask_10_7_7 <= _GEN_2042;
      end
    end else begin
      mask_10_7_7 <= _GEN_2042;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_11_0_0 <= _GEN_8219;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_11_0_0 <= _GEN_4123; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_0 <= 1'h0;
      end else begin
        mask_11_0_0 <= _GEN_1035;
      end
    end else begin
      mask_11_0_0 <= _GEN_1035;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_11_0_1 <= _GEN_8283;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_11_0_1 <= _GEN_4187; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_1 <= 1'h0;
      end else begin
        mask_11_0_1 <= _GEN_1051;
      end
    end else begin
      mask_11_0_1 <= _GEN_1051;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_11_0_2 <= _GEN_8347;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_11_0_2 <= _GEN_4251; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_2 <= 1'h0;
      end else begin
        mask_11_0_2 <= _GEN_1067;
      end
    end else begin
      mask_11_0_2 <= _GEN_1067;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_11_0_3 <= _GEN_8411;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_11_0_3 <= _GEN_4315; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_3 <= 1'h0;
      end else begin
        mask_11_0_3 <= _GEN_1083;
      end
    end else begin
      mask_11_0_3 <= _GEN_1083;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_11_0_4 <= _GEN_8475;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_11_0_4 <= _GEN_4379; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_4 <= 1'h0;
      end else begin
        mask_11_0_4 <= _GEN_1099;
      end
    end else begin
      mask_11_0_4 <= _GEN_1099;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_11_0_5 <= _GEN_8539;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_11_0_5 <= _GEN_4443; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_5 <= 1'h0;
      end else begin
        mask_11_0_5 <= _GEN_1115;
      end
    end else begin
      mask_11_0_5 <= _GEN_1115;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_11_0_6 <= _GEN_8603;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_11_0_6 <= _GEN_4507; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_6 <= 1'h0;
      end else begin
        mask_11_0_6 <= _GEN_1131;
      end
    end else begin
      mask_11_0_6 <= _GEN_1131;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_11_0_7 <= _GEN_8667;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_11_0_7 <= _GEN_4571; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_0_7 <= 1'h0;
      end else begin
        mask_11_0_7 <= _GEN_1147;
      end
    end else begin
      mask_11_0_7 <= _GEN_1147;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_11_1_0 <= _GEN_8731;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_11_1_0 <= _GEN_4635; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_0 <= 1'h0;
      end else begin
        mask_11_1_0 <= _GEN_1163;
      end
    end else begin
      mask_11_1_0 <= _GEN_1163;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_11_1_1 <= _GEN_8795;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_11_1_1 <= _GEN_4699; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_1 <= 1'h0;
      end else begin
        mask_11_1_1 <= _GEN_1179;
      end
    end else begin
      mask_11_1_1 <= _GEN_1179;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_11_1_2 <= _GEN_8859;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_11_1_2 <= _GEN_4763; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_2 <= 1'h0;
      end else begin
        mask_11_1_2 <= _GEN_1195;
      end
    end else begin
      mask_11_1_2 <= _GEN_1195;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_11_1_3 <= _GEN_8923;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_11_1_3 <= _GEN_4827; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_3 <= 1'h0;
      end else begin
        mask_11_1_3 <= _GEN_1211;
      end
    end else begin
      mask_11_1_3 <= _GEN_1211;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_11_1_4 <= _GEN_8987;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_11_1_4 <= _GEN_4891; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_4 <= 1'h0;
      end else begin
        mask_11_1_4 <= _GEN_1227;
      end
    end else begin
      mask_11_1_4 <= _GEN_1227;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_11_1_5 <= _GEN_9051;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_11_1_5 <= _GEN_4955; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_5 <= 1'h0;
      end else begin
        mask_11_1_5 <= _GEN_1243;
      end
    end else begin
      mask_11_1_5 <= _GEN_1243;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_11_1_6 <= _GEN_9115;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_11_1_6 <= _GEN_5019; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_6 <= 1'h0;
      end else begin
        mask_11_1_6 <= _GEN_1259;
      end
    end else begin
      mask_11_1_6 <= _GEN_1259;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_11_1_7 <= _GEN_9179;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_11_1_7 <= _GEN_5083; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_1_7 <= 1'h0;
      end else begin
        mask_11_1_7 <= _GEN_1275;
      end
    end else begin
      mask_11_1_7 <= _GEN_1275;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_11_2_0 <= _GEN_9243;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_11_2_0 <= _GEN_5147; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_0 <= 1'h0;
      end else begin
        mask_11_2_0 <= _GEN_1291;
      end
    end else begin
      mask_11_2_0 <= _GEN_1291;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_11_2_1 <= _GEN_9307;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_11_2_1 <= _GEN_5211; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_1 <= 1'h0;
      end else begin
        mask_11_2_1 <= _GEN_1307;
      end
    end else begin
      mask_11_2_1 <= _GEN_1307;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_11_2_2 <= _GEN_9371;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_11_2_2 <= _GEN_5275; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_2 <= 1'h0;
      end else begin
        mask_11_2_2 <= _GEN_1323;
      end
    end else begin
      mask_11_2_2 <= _GEN_1323;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_11_2_3 <= _GEN_9435;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_11_2_3 <= _GEN_5339; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_3 <= 1'h0;
      end else begin
        mask_11_2_3 <= _GEN_1339;
      end
    end else begin
      mask_11_2_3 <= _GEN_1339;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_11_2_4 <= _GEN_9499;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_11_2_4 <= _GEN_5403; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_4 <= 1'h0;
      end else begin
        mask_11_2_4 <= _GEN_1355;
      end
    end else begin
      mask_11_2_4 <= _GEN_1355;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_11_2_5 <= _GEN_9563;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_11_2_5 <= _GEN_5467; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_5 <= 1'h0;
      end else begin
        mask_11_2_5 <= _GEN_1371;
      end
    end else begin
      mask_11_2_5 <= _GEN_1371;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_11_2_6 <= _GEN_9627;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_11_2_6 <= _GEN_5531; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_6 <= 1'h0;
      end else begin
        mask_11_2_6 <= _GEN_1387;
      end
    end else begin
      mask_11_2_6 <= _GEN_1387;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_11_2_7 <= _GEN_9691;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_11_2_7 <= _GEN_5595; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_2_7 <= 1'h0;
      end else begin
        mask_11_2_7 <= _GEN_1403;
      end
    end else begin
      mask_11_2_7 <= _GEN_1403;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_11_3_0 <= _GEN_9755;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_11_3_0 <= _GEN_5659; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_0 <= 1'h0;
      end else begin
        mask_11_3_0 <= _GEN_1419;
      end
    end else begin
      mask_11_3_0 <= _GEN_1419;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_11_3_1 <= _GEN_9819;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_11_3_1 <= _GEN_5723; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_1 <= 1'h0;
      end else begin
        mask_11_3_1 <= _GEN_1435;
      end
    end else begin
      mask_11_3_1 <= _GEN_1435;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_11_3_2 <= _GEN_9883;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_11_3_2 <= _GEN_5787; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_2 <= 1'h0;
      end else begin
        mask_11_3_2 <= _GEN_1451;
      end
    end else begin
      mask_11_3_2 <= _GEN_1451;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_11_3_3 <= _GEN_9947;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_11_3_3 <= _GEN_5851; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_3 <= 1'h0;
      end else begin
        mask_11_3_3 <= _GEN_1467;
      end
    end else begin
      mask_11_3_3 <= _GEN_1467;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_11_3_4 <= _GEN_10011;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_11_3_4 <= _GEN_5915; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_4 <= 1'h0;
      end else begin
        mask_11_3_4 <= _GEN_1483;
      end
    end else begin
      mask_11_3_4 <= _GEN_1483;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_11_3_5 <= _GEN_10075;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_11_3_5 <= _GEN_5979; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_5 <= 1'h0;
      end else begin
        mask_11_3_5 <= _GEN_1499;
      end
    end else begin
      mask_11_3_5 <= _GEN_1499;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_11_3_6 <= _GEN_10139;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_11_3_6 <= _GEN_6043; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_6 <= 1'h0;
      end else begin
        mask_11_3_6 <= _GEN_1515;
      end
    end else begin
      mask_11_3_6 <= _GEN_1515;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_11_3_7 <= _GEN_10203;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_11_3_7 <= _GEN_6107; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_3_7 <= 1'h0;
      end else begin
        mask_11_3_7 <= _GEN_1531;
      end
    end else begin
      mask_11_3_7 <= _GEN_1531;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_11_4_0 <= _GEN_10267;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_11_4_0 <= _GEN_6171; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_0 <= 1'h0;
      end else begin
        mask_11_4_0 <= _GEN_1547;
      end
    end else begin
      mask_11_4_0 <= _GEN_1547;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_11_4_1 <= _GEN_10331;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_11_4_1 <= _GEN_6235; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_1 <= 1'h0;
      end else begin
        mask_11_4_1 <= _GEN_1563;
      end
    end else begin
      mask_11_4_1 <= _GEN_1563;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_11_4_2 <= _GEN_10395;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_11_4_2 <= _GEN_6299; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_2 <= 1'h0;
      end else begin
        mask_11_4_2 <= _GEN_1579;
      end
    end else begin
      mask_11_4_2 <= _GEN_1579;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_11_4_3 <= _GEN_10459;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_11_4_3 <= _GEN_6363; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_3 <= 1'h0;
      end else begin
        mask_11_4_3 <= _GEN_1595;
      end
    end else begin
      mask_11_4_3 <= _GEN_1595;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_11_4_4 <= _GEN_10523;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_11_4_4 <= _GEN_6427; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_4 <= 1'h0;
      end else begin
        mask_11_4_4 <= _GEN_1611;
      end
    end else begin
      mask_11_4_4 <= _GEN_1611;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_11_4_5 <= _GEN_10587;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_11_4_5 <= _GEN_6491; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_5 <= 1'h0;
      end else begin
        mask_11_4_5 <= _GEN_1627;
      end
    end else begin
      mask_11_4_5 <= _GEN_1627;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_11_4_6 <= _GEN_10651;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_11_4_6 <= _GEN_6555; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_6 <= 1'h0;
      end else begin
        mask_11_4_6 <= _GEN_1643;
      end
    end else begin
      mask_11_4_6 <= _GEN_1643;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_11_4_7 <= _GEN_10715;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_11_4_7 <= _GEN_6619; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_4_7 <= 1'h0;
      end else begin
        mask_11_4_7 <= _GEN_1659;
      end
    end else begin
      mask_11_4_7 <= _GEN_1659;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_11_5_0 <= _GEN_10779;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_11_5_0 <= _GEN_6683; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_0 <= 1'h0;
      end else begin
        mask_11_5_0 <= _GEN_1675;
      end
    end else begin
      mask_11_5_0 <= _GEN_1675;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_11_5_1 <= _GEN_10843;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_11_5_1 <= _GEN_6747; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_1 <= 1'h0;
      end else begin
        mask_11_5_1 <= _GEN_1691;
      end
    end else begin
      mask_11_5_1 <= _GEN_1691;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_11_5_2 <= _GEN_10907;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_11_5_2 <= _GEN_6811; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_2 <= 1'h0;
      end else begin
        mask_11_5_2 <= _GEN_1707;
      end
    end else begin
      mask_11_5_2 <= _GEN_1707;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_11_5_3 <= _GEN_10971;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_11_5_3 <= _GEN_6875; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_3 <= 1'h0;
      end else begin
        mask_11_5_3 <= _GEN_1723;
      end
    end else begin
      mask_11_5_3 <= _GEN_1723;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_11_5_4 <= _GEN_11035;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_11_5_4 <= _GEN_6939; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_4 <= 1'h0;
      end else begin
        mask_11_5_4 <= _GEN_1739;
      end
    end else begin
      mask_11_5_4 <= _GEN_1739;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_11_5_5 <= _GEN_11099;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_11_5_5 <= _GEN_7003; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_5 <= 1'h0;
      end else begin
        mask_11_5_5 <= _GEN_1755;
      end
    end else begin
      mask_11_5_5 <= _GEN_1755;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_11_5_6 <= _GEN_11163;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_11_5_6 <= _GEN_7067; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_6 <= 1'h0;
      end else begin
        mask_11_5_6 <= _GEN_1771;
      end
    end else begin
      mask_11_5_6 <= _GEN_1771;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_11_5_7 <= _GEN_11227;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_11_5_7 <= _GEN_7131; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_5_7 <= 1'h0;
      end else begin
        mask_11_5_7 <= _GEN_1787;
      end
    end else begin
      mask_11_5_7 <= _GEN_1787;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_11_6_0 <= _GEN_11291;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_11_6_0 <= _GEN_7195; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_0 <= 1'h0;
      end else begin
        mask_11_6_0 <= _GEN_1803;
      end
    end else begin
      mask_11_6_0 <= _GEN_1803;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_11_6_1 <= _GEN_11355;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_11_6_1 <= _GEN_7259; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_1 <= 1'h0;
      end else begin
        mask_11_6_1 <= _GEN_1819;
      end
    end else begin
      mask_11_6_1 <= _GEN_1819;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_11_6_2 <= _GEN_11419;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_11_6_2 <= _GEN_7323; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_2 <= 1'h0;
      end else begin
        mask_11_6_2 <= _GEN_1835;
      end
    end else begin
      mask_11_6_2 <= _GEN_1835;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_11_6_3 <= _GEN_11483;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_11_6_3 <= _GEN_7387; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_3 <= 1'h0;
      end else begin
        mask_11_6_3 <= _GEN_1851;
      end
    end else begin
      mask_11_6_3 <= _GEN_1851;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_11_6_4 <= _GEN_11547;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_11_6_4 <= _GEN_7451; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_4 <= 1'h0;
      end else begin
        mask_11_6_4 <= _GEN_1867;
      end
    end else begin
      mask_11_6_4 <= _GEN_1867;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_11_6_5 <= _GEN_11611;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_11_6_5 <= _GEN_7515; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_5 <= 1'h0;
      end else begin
        mask_11_6_5 <= _GEN_1883;
      end
    end else begin
      mask_11_6_5 <= _GEN_1883;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_11_6_6 <= _GEN_11675;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_11_6_6 <= _GEN_7579; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_6 <= 1'h0;
      end else begin
        mask_11_6_6 <= _GEN_1899;
      end
    end else begin
      mask_11_6_6 <= _GEN_1899;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_11_6_7 <= _GEN_11739;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_11_6_7 <= _GEN_7643; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_6_7 <= 1'h0;
      end else begin
        mask_11_6_7 <= _GEN_1915;
      end
    end else begin
      mask_11_6_7 <= _GEN_1915;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_11_7_0 <= _GEN_11803;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_11_7_0 <= _GEN_7707; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_0 <= 1'h0;
      end else begin
        mask_11_7_0 <= _GEN_1931;
      end
    end else begin
      mask_11_7_0 <= _GEN_1931;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_11_7_1 <= _GEN_11867;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_11_7_1 <= _GEN_7771; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_1 <= 1'h0;
      end else begin
        mask_11_7_1 <= _GEN_1947;
      end
    end else begin
      mask_11_7_1 <= _GEN_1947;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_11_7_2 <= _GEN_11931;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_11_7_2 <= _GEN_7835; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_2 <= 1'h0;
      end else begin
        mask_11_7_2 <= _GEN_1963;
      end
    end else begin
      mask_11_7_2 <= _GEN_1963;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_11_7_3 <= _GEN_11995;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_11_7_3 <= _GEN_7899; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_3 <= 1'h0;
      end else begin
        mask_11_7_3 <= _GEN_1979;
      end
    end else begin
      mask_11_7_3 <= _GEN_1979;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_11_7_4 <= _GEN_12059;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_11_7_4 <= _GEN_7963; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_4 <= 1'h0;
      end else begin
        mask_11_7_4 <= _GEN_1995;
      end
    end else begin
      mask_11_7_4 <= _GEN_1995;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_11_7_5 <= _GEN_12123;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_11_7_5 <= _GEN_8027; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_5 <= 1'h0;
      end else begin
        mask_11_7_5 <= _GEN_2011;
      end
    end else begin
      mask_11_7_5 <= _GEN_2011;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_11_7_6 <= _GEN_12187;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_11_7_6 <= _GEN_8091; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_6 <= 1'h0;
      end else begin
        mask_11_7_6 <= _GEN_2027;
      end
    end else begin
      mask_11_7_6 <= _GEN_2027;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_11_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_11_7_7 <= _GEN_12251;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_11_7_7 <= _GEN_8155; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hb == line_mask_clean_line_1) begin
        mask_11_7_7 <= 1'h0;
      end else begin
        mask_11_7_7 <= _GEN_2043;
      end
    end else begin
      mask_11_7_7 <= _GEN_2043;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_12_0_0 <= _GEN_8220;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_12_0_0 <= _GEN_4124; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_0 <= 1'h0;
      end else begin
        mask_12_0_0 <= _GEN_1036;
      end
    end else begin
      mask_12_0_0 <= _GEN_1036;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_12_0_1 <= _GEN_8284;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_12_0_1 <= _GEN_4188; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_1 <= 1'h0;
      end else begin
        mask_12_0_1 <= _GEN_1052;
      end
    end else begin
      mask_12_0_1 <= _GEN_1052;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_12_0_2 <= _GEN_8348;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_12_0_2 <= _GEN_4252; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_2 <= 1'h0;
      end else begin
        mask_12_0_2 <= _GEN_1068;
      end
    end else begin
      mask_12_0_2 <= _GEN_1068;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_12_0_3 <= _GEN_8412;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_12_0_3 <= _GEN_4316; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_3 <= 1'h0;
      end else begin
        mask_12_0_3 <= _GEN_1084;
      end
    end else begin
      mask_12_0_3 <= _GEN_1084;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_12_0_4 <= _GEN_8476;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_12_0_4 <= _GEN_4380; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_4 <= 1'h0;
      end else begin
        mask_12_0_4 <= _GEN_1100;
      end
    end else begin
      mask_12_0_4 <= _GEN_1100;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_12_0_5 <= _GEN_8540;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_12_0_5 <= _GEN_4444; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_5 <= 1'h0;
      end else begin
        mask_12_0_5 <= _GEN_1116;
      end
    end else begin
      mask_12_0_5 <= _GEN_1116;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_12_0_6 <= _GEN_8604;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_12_0_6 <= _GEN_4508; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_6 <= 1'h0;
      end else begin
        mask_12_0_6 <= _GEN_1132;
      end
    end else begin
      mask_12_0_6 <= _GEN_1132;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_12_0_7 <= _GEN_8668;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_12_0_7 <= _GEN_4572; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_0_7 <= 1'h0;
      end else begin
        mask_12_0_7 <= _GEN_1148;
      end
    end else begin
      mask_12_0_7 <= _GEN_1148;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_12_1_0 <= _GEN_8732;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_12_1_0 <= _GEN_4636; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_0 <= 1'h0;
      end else begin
        mask_12_1_0 <= _GEN_1164;
      end
    end else begin
      mask_12_1_0 <= _GEN_1164;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_12_1_1 <= _GEN_8796;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_12_1_1 <= _GEN_4700; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_1 <= 1'h0;
      end else begin
        mask_12_1_1 <= _GEN_1180;
      end
    end else begin
      mask_12_1_1 <= _GEN_1180;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_12_1_2 <= _GEN_8860;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_12_1_2 <= _GEN_4764; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_2 <= 1'h0;
      end else begin
        mask_12_1_2 <= _GEN_1196;
      end
    end else begin
      mask_12_1_2 <= _GEN_1196;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_12_1_3 <= _GEN_8924;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_12_1_3 <= _GEN_4828; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_3 <= 1'h0;
      end else begin
        mask_12_1_3 <= _GEN_1212;
      end
    end else begin
      mask_12_1_3 <= _GEN_1212;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_12_1_4 <= _GEN_8988;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_12_1_4 <= _GEN_4892; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_4 <= 1'h0;
      end else begin
        mask_12_1_4 <= _GEN_1228;
      end
    end else begin
      mask_12_1_4 <= _GEN_1228;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_12_1_5 <= _GEN_9052;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_12_1_5 <= _GEN_4956; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_5 <= 1'h0;
      end else begin
        mask_12_1_5 <= _GEN_1244;
      end
    end else begin
      mask_12_1_5 <= _GEN_1244;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_12_1_6 <= _GEN_9116;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_12_1_6 <= _GEN_5020; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_6 <= 1'h0;
      end else begin
        mask_12_1_6 <= _GEN_1260;
      end
    end else begin
      mask_12_1_6 <= _GEN_1260;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_12_1_7 <= _GEN_9180;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_12_1_7 <= _GEN_5084; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_1_7 <= 1'h0;
      end else begin
        mask_12_1_7 <= _GEN_1276;
      end
    end else begin
      mask_12_1_7 <= _GEN_1276;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_12_2_0 <= _GEN_9244;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_12_2_0 <= _GEN_5148; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_0 <= 1'h0;
      end else begin
        mask_12_2_0 <= _GEN_1292;
      end
    end else begin
      mask_12_2_0 <= _GEN_1292;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_12_2_1 <= _GEN_9308;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_12_2_1 <= _GEN_5212; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_1 <= 1'h0;
      end else begin
        mask_12_2_1 <= _GEN_1308;
      end
    end else begin
      mask_12_2_1 <= _GEN_1308;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_12_2_2 <= _GEN_9372;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_12_2_2 <= _GEN_5276; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_2 <= 1'h0;
      end else begin
        mask_12_2_2 <= _GEN_1324;
      end
    end else begin
      mask_12_2_2 <= _GEN_1324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_12_2_3 <= _GEN_9436;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_12_2_3 <= _GEN_5340; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_3 <= 1'h0;
      end else begin
        mask_12_2_3 <= _GEN_1340;
      end
    end else begin
      mask_12_2_3 <= _GEN_1340;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_12_2_4 <= _GEN_9500;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_12_2_4 <= _GEN_5404; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_4 <= 1'h0;
      end else begin
        mask_12_2_4 <= _GEN_1356;
      end
    end else begin
      mask_12_2_4 <= _GEN_1356;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_12_2_5 <= _GEN_9564;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_12_2_5 <= _GEN_5468; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_5 <= 1'h0;
      end else begin
        mask_12_2_5 <= _GEN_1372;
      end
    end else begin
      mask_12_2_5 <= _GEN_1372;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_12_2_6 <= _GEN_9628;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_12_2_6 <= _GEN_5532; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_6 <= 1'h0;
      end else begin
        mask_12_2_6 <= _GEN_1388;
      end
    end else begin
      mask_12_2_6 <= _GEN_1388;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_12_2_7 <= _GEN_9692;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_12_2_7 <= _GEN_5596; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_2_7 <= 1'h0;
      end else begin
        mask_12_2_7 <= _GEN_1404;
      end
    end else begin
      mask_12_2_7 <= _GEN_1404;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_12_3_0 <= _GEN_9756;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_12_3_0 <= _GEN_5660; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_0 <= 1'h0;
      end else begin
        mask_12_3_0 <= _GEN_1420;
      end
    end else begin
      mask_12_3_0 <= _GEN_1420;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_12_3_1 <= _GEN_9820;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_12_3_1 <= _GEN_5724; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_1 <= 1'h0;
      end else begin
        mask_12_3_1 <= _GEN_1436;
      end
    end else begin
      mask_12_3_1 <= _GEN_1436;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_12_3_2 <= _GEN_9884;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_12_3_2 <= _GEN_5788; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_2 <= 1'h0;
      end else begin
        mask_12_3_2 <= _GEN_1452;
      end
    end else begin
      mask_12_3_2 <= _GEN_1452;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_12_3_3 <= _GEN_9948;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_12_3_3 <= _GEN_5852; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_3 <= 1'h0;
      end else begin
        mask_12_3_3 <= _GEN_1468;
      end
    end else begin
      mask_12_3_3 <= _GEN_1468;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_12_3_4 <= _GEN_10012;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_12_3_4 <= _GEN_5916; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_4 <= 1'h0;
      end else begin
        mask_12_3_4 <= _GEN_1484;
      end
    end else begin
      mask_12_3_4 <= _GEN_1484;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_12_3_5 <= _GEN_10076;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_12_3_5 <= _GEN_5980; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_5 <= 1'h0;
      end else begin
        mask_12_3_5 <= _GEN_1500;
      end
    end else begin
      mask_12_3_5 <= _GEN_1500;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_12_3_6 <= _GEN_10140;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_12_3_6 <= _GEN_6044; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_6 <= 1'h0;
      end else begin
        mask_12_3_6 <= _GEN_1516;
      end
    end else begin
      mask_12_3_6 <= _GEN_1516;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_12_3_7 <= _GEN_10204;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_12_3_7 <= _GEN_6108; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_3_7 <= 1'h0;
      end else begin
        mask_12_3_7 <= _GEN_1532;
      end
    end else begin
      mask_12_3_7 <= _GEN_1532;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_12_4_0 <= _GEN_10268;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_12_4_0 <= _GEN_6172; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_0 <= 1'h0;
      end else begin
        mask_12_4_0 <= _GEN_1548;
      end
    end else begin
      mask_12_4_0 <= _GEN_1548;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_12_4_1 <= _GEN_10332;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_12_4_1 <= _GEN_6236; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_1 <= 1'h0;
      end else begin
        mask_12_4_1 <= _GEN_1564;
      end
    end else begin
      mask_12_4_1 <= _GEN_1564;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_12_4_2 <= _GEN_10396;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_12_4_2 <= _GEN_6300; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_2 <= 1'h0;
      end else begin
        mask_12_4_2 <= _GEN_1580;
      end
    end else begin
      mask_12_4_2 <= _GEN_1580;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_12_4_3 <= _GEN_10460;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_12_4_3 <= _GEN_6364; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_3 <= 1'h0;
      end else begin
        mask_12_4_3 <= _GEN_1596;
      end
    end else begin
      mask_12_4_3 <= _GEN_1596;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_12_4_4 <= _GEN_10524;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_12_4_4 <= _GEN_6428; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_4 <= 1'h0;
      end else begin
        mask_12_4_4 <= _GEN_1612;
      end
    end else begin
      mask_12_4_4 <= _GEN_1612;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_12_4_5 <= _GEN_10588;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_12_4_5 <= _GEN_6492; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_5 <= 1'h0;
      end else begin
        mask_12_4_5 <= _GEN_1628;
      end
    end else begin
      mask_12_4_5 <= _GEN_1628;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_12_4_6 <= _GEN_10652;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_12_4_6 <= _GEN_6556; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_6 <= 1'h0;
      end else begin
        mask_12_4_6 <= _GEN_1644;
      end
    end else begin
      mask_12_4_6 <= _GEN_1644;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_12_4_7 <= _GEN_10716;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_12_4_7 <= _GEN_6620; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_4_7 <= 1'h0;
      end else begin
        mask_12_4_7 <= _GEN_1660;
      end
    end else begin
      mask_12_4_7 <= _GEN_1660;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_12_5_0 <= _GEN_10780;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_12_5_0 <= _GEN_6684; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_0 <= 1'h0;
      end else begin
        mask_12_5_0 <= _GEN_1676;
      end
    end else begin
      mask_12_5_0 <= _GEN_1676;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_12_5_1 <= _GEN_10844;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_12_5_1 <= _GEN_6748; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_1 <= 1'h0;
      end else begin
        mask_12_5_1 <= _GEN_1692;
      end
    end else begin
      mask_12_5_1 <= _GEN_1692;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_12_5_2 <= _GEN_10908;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_12_5_2 <= _GEN_6812; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_2 <= 1'h0;
      end else begin
        mask_12_5_2 <= _GEN_1708;
      end
    end else begin
      mask_12_5_2 <= _GEN_1708;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_12_5_3 <= _GEN_10972;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_12_5_3 <= _GEN_6876; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_3 <= 1'h0;
      end else begin
        mask_12_5_3 <= _GEN_1724;
      end
    end else begin
      mask_12_5_3 <= _GEN_1724;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_12_5_4 <= _GEN_11036;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_12_5_4 <= _GEN_6940; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_4 <= 1'h0;
      end else begin
        mask_12_5_4 <= _GEN_1740;
      end
    end else begin
      mask_12_5_4 <= _GEN_1740;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_12_5_5 <= _GEN_11100;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_12_5_5 <= _GEN_7004; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_5 <= 1'h0;
      end else begin
        mask_12_5_5 <= _GEN_1756;
      end
    end else begin
      mask_12_5_5 <= _GEN_1756;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_12_5_6 <= _GEN_11164;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_12_5_6 <= _GEN_7068; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_6 <= 1'h0;
      end else begin
        mask_12_5_6 <= _GEN_1772;
      end
    end else begin
      mask_12_5_6 <= _GEN_1772;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_12_5_7 <= _GEN_11228;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_12_5_7 <= _GEN_7132; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_5_7 <= 1'h0;
      end else begin
        mask_12_5_7 <= _GEN_1788;
      end
    end else begin
      mask_12_5_7 <= _GEN_1788;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_12_6_0 <= _GEN_11292;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_12_6_0 <= _GEN_7196; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_0 <= 1'h0;
      end else begin
        mask_12_6_0 <= _GEN_1804;
      end
    end else begin
      mask_12_6_0 <= _GEN_1804;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_12_6_1 <= _GEN_11356;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_12_6_1 <= _GEN_7260; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_1 <= 1'h0;
      end else begin
        mask_12_6_1 <= _GEN_1820;
      end
    end else begin
      mask_12_6_1 <= _GEN_1820;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_12_6_2 <= _GEN_11420;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_12_6_2 <= _GEN_7324; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_2 <= 1'h0;
      end else begin
        mask_12_6_2 <= _GEN_1836;
      end
    end else begin
      mask_12_6_2 <= _GEN_1836;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_12_6_3 <= _GEN_11484;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_12_6_3 <= _GEN_7388; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_3 <= 1'h0;
      end else begin
        mask_12_6_3 <= _GEN_1852;
      end
    end else begin
      mask_12_6_3 <= _GEN_1852;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_12_6_4 <= _GEN_11548;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_12_6_4 <= _GEN_7452; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_4 <= 1'h0;
      end else begin
        mask_12_6_4 <= _GEN_1868;
      end
    end else begin
      mask_12_6_4 <= _GEN_1868;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_12_6_5 <= _GEN_11612;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_12_6_5 <= _GEN_7516; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_5 <= 1'h0;
      end else begin
        mask_12_6_5 <= _GEN_1884;
      end
    end else begin
      mask_12_6_5 <= _GEN_1884;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_12_6_6 <= _GEN_11676;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_12_6_6 <= _GEN_7580; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_6 <= 1'h0;
      end else begin
        mask_12_6_6 <= _GEN_1900;
      end
    end else begin
      mask_12_6_6 <= _GEN_1900;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_12_6_7 <= _GEN_11740;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_12_6_7 <= _GEN_7644; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_6_7 <= 1'h0;
      end else begin
        mask_12_6_7 <= _GEN_1916;
      end
    end else begin
      mask_12_6_7 <= _GEN_1916;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_12_7_0 <= _GEN_11804;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_12_7_0 <= _GEN_7708; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_0 <= 1'h0;
      end else begin
        mask_12_7_0 <= _GEN_1932;
      end
    end else begin
      mask_12_7_0 <= _GEN_1932;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_12_7_1 <= _GEN_11868;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_12_7_1 <= _GEN_7772; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_1 <= 1'h0;
      end else begin
        mask_12_7_1 <= _GEN_1948;
      end
    end else begin
      mask_12_7_1 <= _GEN_1948;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_12_7_2 <= _GEN_11932;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_12_7_2 <= _GEN_7836; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_2 <= 1'h0;
      end else begin
        mask_12_7_2 <= _GEN_1964;
      end
    end else begin
      mask_12_7_2 <= _GEN_1964;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_12_7_3 <= _GEN_11996;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_12_7_3 <= _GEN_7900; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_3 <= 1'h0;
      end else begin
        mask_12_7_3 <= _GEN_1980;
      end
    end else begin
      mask_12_7_3 <= _GEN_1980;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_12_7_4 <= _GEN_12060;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_12_7_4 <= _GEN_7964; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_4 <= 1'h0;
      end else begin
        mask_12_7_4 <= _GEN_1996;
      end
    end else begin
      mask_12_7_4 <= _GEN_1996;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_12_7_5 <= _GEN_12124;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_12_7_5 <= _GEN_8028; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_5 <= 1'h0;
      end else begin
        mask_12_7_5 <= _GEN_2012;
      end
    end else begin
      mask_12_7_5 <= _GEN_2012;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_12_7_6 <= _GEN_12188;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_12_7_6 <= _GEN_8092; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_6 <= 1'h0;
      end else begin
        mask_12_7_6 <= _GEN_2028;
      end
    end else begin
      mask_12_7_6 <= _GEN_2028;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_12_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_12_7_7 <= _GEN_12252;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_12_7_7 <= _GEN_8156; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hc == line_mask_clean_line_1) begin
        mask_12_7_7 <= 1'h0;
      end else begin
        mask_12_7_7 <= _GEN_2044;
      end
    end else begin
      mask_12_7_7 <= _GEN_2044;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_13_0_0 <= _GEN_8221;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_13_0_0 <= _GEN_4125; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_0 <= 1'h0;
      end else begin
        mask_13_0_0 <= _GEN_1037;
      end
    end else begin
      mask_13_0_0 <= _GEN_1037;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_13_0_1 <= _GEN_8285;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_13_0_1 <= _GEN_4189; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_1 <= 1'h0;
      end else begin
        mask_13_0_1 <= _GEN_1053;
      end
    end else begin
      mask_13_0_1 <= _GEN_1053;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_13_0_2 <= _GEN_8349;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_13_0_2 <= _GEN_4253; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_2 <= 1'h0;
      end else begin
        mask_13_0_2 <= _GEN_1069;
      end
    end else begin
      mask_13_0_2 <= _GEN_1069;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_13_0_3 <= _GEN_8413;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_13_0_3 <= _GEN_4317; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_3 <= 1'h0;
      end else begin
        mask_13_0_3 <= _GEN_1085;
      end
    end else begin
      mask_13_0_3 <= _GEN_1085;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_13_0_4 <= _GEN_8477;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_13_0_4 <= _GEN_4381; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_4 <= 1'h0;
      end else begin
        mask_13_0_4 <= _GEN_1101;
      end
    end else begin
      mask_13_0_4 <= _GEN_1101;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_13_0_5 <= _GEN_8541;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_13_0_5 <= _GEN_4445; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_5 <= 1'h0;
      end else begin
        mask_13_0_5 <= _GEN_1117;
      end
    end else begin
      mask_13_0_5 <= _GEN_1117;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_13_0_6 <= _GEN_8605;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_13_0_6 <= _GEN_4509; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_6 <= 1'h0;
      end else begin
        mask_13_0_6 <= _GEN_1133;
      end
    end else begin
      mask_13_0_6 <= _GEN_1133;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_13_0_7 <= _GEN_8669;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_13_0_7 <= _GEN_4573; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_0_7 <= 1'h0;
      end else begin
        mask_13_0_7 <= _GEN_1149;
      end
    end else begin
      mask_13_0_7 <= _GEN_1149;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_13_1_0 <= _GEN_8733;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_13_1_0 <= _GEN_4637; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_0 <= 1'h0;
      end else begin
        mask_13_1_0 <= _GEN_1165;
      end
    end else begin
      mask_13_1_0 <= _GEN_1165;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_13_1_1 <= _GEN_8797;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_13_1_1 <= _GEN_4701; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_1 <= 1'h0;
      end else begin
        mask_13_1_1 <= _GEN_1181;
      end
    end else begin
      mask_13_1_1 <= _GEN_1181;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_13_1_2 <= _GEN_8861;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_13_1_2 <= _GEN_4765; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_2 <= 1'h0;
      end else begin
        mask_13_1_2 <= _GEN_1197;
      end
    end else begin
      mask_13_1_2 <= _GEN_1197;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_13_1_3 <= _GEN_8925;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_13_1_3 <= _GEN_4829; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_3 <= 1'h0;
      end else begin
        mask_13_1_3 <= _GEN_1213;
      end
    end else begin
      mask_13_1_3 <= _GEN_1213;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_13_1_4 <= _GEN_8989;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_13_1_4 <= _GEN_4893; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_4 <= 1'h0;
      end else begin
        mask_13_1_4 <= _GEN_1229;
      end
    end else begin
      mask_13_1_4 <= _GEN_1229;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_13_1_5 <= _GEN_9053;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_13_1_5 <= _GEN_4957; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_5 <= 1'h0;
      end else begin
        mask_13_1_5 <= _GEN_1245;
      end
    end else begin
      mask_13_1_5 <= _GEN_1245;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_13_1_6 <= _GEN_9117;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_13_1_6 <= _GEN_5021; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_6 <= 1'h0;
      end else begin
        mask_13_1_6 <= _GEN_1261;
      end
    end else begin
      mask_13_1_6 <= _GEN_1261;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_13_1_7 <= _GEN_9181;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_13_1_7 <= _GEN_5085; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_1_7 <= 1'h0;
      end else begin
        mask_13_1_7 <= _GEN_1277;
      end
    end else begin
      mask_13_1_7 <= _GEN_1277;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_13_2_0 <= _GEN_9245;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_13_2_0 <= _GEN_5149; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_0 <= 1'h0;
      end else begin
        mask_13_2_0 <= _GEN_1293;
      end
    end else begin
      mask_13_2_0 <= _GEN_1293;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_13_2_1 <= _GEN_9309;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_13_2_1 <= _GEN_5213; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_1 <= 1'h0;
      end else begin
        mask_13_2_1 <= _GEN_1309;
      end
    end else begin
      mask_13_2_1 <= _GEN_1309;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_13_2_2 <= _GEN_9373;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_13_2_2 <= _GEN_5277; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_2 <= 1'h0;
      end else begin
        mask_13_2_2 <= _GEN_1325;
      end
    end else begin
      mask_13_2_2 <= _GEN_1325;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_13_2_3 <= _GEN_9437;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_13_2_3 <= _GEN_5341; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_3 <= 1'h0;
      end else begin
        mask_13_2_3 <= _GEN_1341;
      end
    end else begin
      mask_13_2_3 <= _GEN_1341;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_13_2_4 <= _GEN_9501;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_13_2_4 <= _GEN_5405; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_4 <= 1'h0;
      end else begin
        mask_13_2_4 <= _GEN_1357;
      end
    end else begin
      mask_13_2_4 <= _GEN_1357;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_13_2_5 <= _GEN_9565;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_13_2_5 <= _GEN_5469; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_5 <= 1'h0;
      end else begin
        mask_13_2_5 <= _GEN_1373;
      end
    end else begin
      mask_13_2_5 <= _GEN_1373;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_13_2_6 <= _GEN_9629;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_13_2_6 <= _GEN_5533; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_6 <= 1'h0;
      end else begin
        mask_13_2_6 <= _GEN_1389;
      end
    end else begin
      mask_13_2_6 <= _GEN_1389;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_13_2_7 <= _GEN_9693;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_13_2_7 <= _GEN_5597; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_2_7 <= 1'h0;
      end else begin
        mask_13_2_7 <= _GEN_1405;
      end
    end else begin
      mask_13_2_7 <= _GEN_1405;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_13_3_0 <= _GEN_9757;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_13_3_0 <= _GEN_5661; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_0 <= 1'h0;
      end else begin
        mask_13_3_0 <= _GEN_1421;
      end
    end else begin
      mask_13_3_0 <= _GEN_1421;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_13_3_1 <= _GEN_9821;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_13_3_1 <= _GEN_5725; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_1 <= 1'h0;
      end else begin
        mask_13_3_1 <= _GEN_1437;
      end
    end else begin
      mask_13_3_1 <= _GEN_1437;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_13_3_2 <= _GEN_9885;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_13_3_2 <= _GEN_5789; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_2 <= 1'h0;
      end else begin
        mask_13_3_2 <= _GEN_1453;
      end
    end else begin
      mask_13_3_2 <= _GEN_1453;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_13_3_3 <= _GEN_9949;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_13_3_3 <= _GEN_5853; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_3 <= 1'h0;
      end else begin
        mask_13_3_3 <= _GEN_1469;
      end
    end else begin
      mask_13_3_3 <= _GEN_1469;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_13_3_4 <= _GEN_10013;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_13_3_4 <= _GEN_5917; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_4 <= 1'h0;
      end else begin
        mask_13_3_4 <= _GEN_1485;
      end
    end else begin
      mask_13_3_4 <= _GEN_1485;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_13_3_5 <= _GEN_10077;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_13_3_5 <= _GEN_5981; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_5 <= 1'h0;
      end else begin
        mask_13_3_5 <= _GEN_1501;
      end
    end else begin
      mask_13_3_5 <= _GEN_1501;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_13_3_6 <= _GEN_10141;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_13_3_6 <= _GEN_6045; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_6 <= 1'h0;
      end else begin
        mask_13_3_6 <= _GEN_1517;
      end
    end else begin
      mask_13_3_6 <= _GEN_1517;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_13_3_7 <= _GEN_10205;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_13_3_7 <= _GEN_6109; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_3_7 <= 1'h0;
      end else begin
        mask_13_3_7 <= _GEN_1533;
      end
    end else begin
      mask_13_3_7 <= _GEN_1533;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_13_4_0 <= _GEN_10269;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_13_4_0 <= _GEN_6173; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_0 <= 1'h0;
      end else begin
        mask_13_4_0 <= _GEN_1549;
      end
    end else begin
      mask_13_4_0 <= _GEN_1549;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_13_4_1 <= _GEN_10333;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_13_4_1 <= _GEN_6237; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_1 <= 1'h0;
      end else begin
        mask_13_4_1 <= _GEN_1565;
      end
    end else begin
      mask_13_4_1 <= _GEN_1565;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_13_4_2 <= _GEN_10397;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_13_4_2 <= _GEN_6301; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_2 <= 1'h0;
      end else begin
        mask_13_4_2 <= _GEN_1581;
      end
    end else begin
      mask_13_4_2 <= _GEN_1581;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_13_4_3 <= _GEN_10461;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_13_4_3 <= _GEN_6365; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_3 <= 1'h0;
      end else begin
        mask_13_4_3 <= _GEN_1597;
      end
    end else begin
      mask_13_4_3 <= _GEN_1597;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_13_4_4 <= _GEN_10525;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_13_4_4 <= _GEN_6429; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_4 <= 1'h0;
      end else begin
        mask_13_4_4 <= _GEN_1613;
      end
    end else begin
      mask_13_4_4 <= _GEN_1613;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_13_4_5 <= _GEN_10589;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_13_4_5 <= _GEN_6493; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_5 <= 1'h0;
      end else begin
        mask_13_4_5 <= _GEN_1629;
      end
    end else begin
      mask_13_4_5 <= _GEN_1629;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_13_4_6 <= _GEN_10653;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_13_4_6 <= _GEN_6557; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_6 <= 1'h0;
      end else begin
        mask_13_4_6 <= _GEN_1645;
      end
    end else begin
      mask_13_4_6 <= _GEN_1645;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_13_4_7 <= _GEN_10717;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_13_4_7 <= _GEN_6621; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_4_7 <= 1'h0;
      end else begin
        mask_13_4_7 <= _GEN_1661;
      end
    end else begin
      mask_13_4_7 <= _GEN_1661;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_13_5_0 <= _GEN_10781;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_13_5_0 <= _GEN_6685; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_0 <= 1'h0;
      end else begin
        mask_13_5_0 <= _GEN_1677;
      end
    end else begin
      mask_13_5_0 <= _GEN_1677;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_13_5_1 <= _GEN_10845;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_13_5_1 <= _GEN_6749; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_1 <= 1'h0;
      end else begin
        mask_13_5_1 <= _GEN_1693;
      end
    end else begin
      mask_13_5_1 <= _GEN_1693;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_13_5_2 <= _GEN_10909;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_13_5_2 <= _GEN_6813; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_2 <= 1'h0;
      end else begin
        mask_13_5_2 <= _GEN_1709;
      end
    end else begin
      mask_13_5_2 <= _GEN_1709;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_13_5_3 <= _GEN_10973;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_13_5_3 <= _GEN_6877; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_3 <= 1'h0;
      end else begin
        mask_13_5_3 <= _GEN_1725;
      end
    end else begin
      mask_13_5_3 <= _GEN_1725;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_13_5_4 <= _GEN_11037;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_13_5_4 <= _GEN_6941; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_4 <= 1'h0;
      end else begin
        mask_13_5_4 <= _GEN_1741;
      end
    end else begin
      mask_13_5_4 <= _GEN_1741;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_13_5_5 <= _GEN_11101;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_13_5_5 <= _GEN_7005; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_5 <= 1'h0;
      end else begin
        mask_13_5_5 <= _GEN_1757;
      end
    end else begin
      mask_13_5_5 <= _GEN_1757;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_13_5_6 <= _GEN_11165;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_13_5_6 <= _GEN_7069; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_6 <= 1'h0;
      end else begin
        mask_13_5_6 <= _GEN_1773;
      end
    end else begin
      mask_13_5_6 <= _GEN_1773;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_13_5_7 <= _GEN_11229;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_13_5_7 <= _GEN_7133; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_5_7 <= 1'h0;
      end else begin
        mask_13_5_7 <= _GEN_1789;
      end
    end else begin
      mask_13_5_7 <= _GEN_1789;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_13_6_0 <= _GEN_11293;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_13_6_0 <= _GEN_7197; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_0 <= 1'h0;
      end else begin
        mask_13_6_0 <= _GEN_1805;
      end
    end else begin
      mask_13_6_0 <= _GEN_1805;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_13_6_1 <= _GEN_11357;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_13_6_1 <= _GEN_7261; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_1 <= 1'h0;
      end else begin
        mask_13_6_1 <= _GEN_1821;
      end
    end else begin
      mask_13_6_1 <= _GEN_1821;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_13_6_2 <= _GEN_11421;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_13_6_2 <= _GEN_7325; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_2 <= 1'h0;
      end else begin
        mask_13_6_2 <= _GEN_1837;
      end
    end else begin
      mask_13_6_2 <= _GEN_1837;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_13_6_3 <= _GEN_11485;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_13_6_3 <= _GEN_7389; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_3 <= 1'h0;
      end else begin
        mask_13_6_3 <= _GEN_1853;
      end
    end else begin
      mask_13_6_3 <= _GEN_1853;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_13_6_4 <= _GEN_11549;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_13_6_4 <= _GEN_7453; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_4 <= 1'h0;
      end else begin
        mask_13_6_4 <= _GEN_1869;
      end
    end else begin
      mask_13_6_4 <= _GEN_1869;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_13_6_5 <= _GEN_11613;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_13_6_5 <= _GEN_7517; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_5 <= 1'h0;
      end else begin
        mask_13_6_5 <= _GEN_1885;
      end
    end else begin
      mask_13_6_5 <= _GEN_1885;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_13_6_6 <= _GEN_11677;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_13_6_6 <= _GEN_7581; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_6 <= 1'h0;
      end else begin
        mask_13_6_6 <= _GEN_1901;
      end
    end else begin
      mask_13_6_6 <= _GEN_1901;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_13_6_7 <= _GEN_11741;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_13_6_7 <= _GEN_7645; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_6_7 <= 1'h0;
      end else begin
        mask_13_6_7 <= _GEN_1917;
      end
    end else begin
      mask_13_6_7 <= _GEN_1917;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_13_7_0 <= _GEN_11805;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_13_7_0 <= _GEN_7709; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_0 <= 1'h0;
      end else begin
        mask_13_7_0 <= _GEN_1933;
      end
    end else begin
      mask_13_7_0 <= _GEN_1933;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_13_7_1 <= _GEN_11869;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_13_7_1 <= _GEN_7773; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_1 <= 1'h0;
      end else begin
        mask_13_7_1 <= _GEN_1949;
      end
    end else begin
      mask_13_7_1 <= _GEN_1949;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_13_7_2 <= _GEN_11933;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_13_7_2 <= _GEN_7837; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_2 <= 1'h0;
      end else begin
        mask_13_7_2 <= _GEN_1965;
      end
    end else begin
      mask_13_7_2 <= _GEN_1965;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_13_7_3 <= _GEN_11997;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_13_7_3 <= _GEN_7901; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_3 <= 1'h0;
      end else begin
        mask_13_7_3 <= _GEN_1981;
      end
    end else begin
      mask_13_7_3 <= _GEN_1981;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_13_7_4 <= _GEN_12061;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_13_7_4 <= _GEN_7965; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_4 <= 1'h0;
      end else begin
        mask_13_7_4 <= _GEN_1997;
      end
    end else begin
      mask_13_7_4 <= _GEN_1997;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_13_7_5 <= _GEN_12125;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_13_7_5 <= _GEN_8029; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_5 <= 1'h0;
      end else begin
        mask_13_7_5 <= _GEN_2013;
      end
    end else begin
      mask_13_7_5 <= _GEN_2013;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_13_7_6 <= _GEN_12189;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_13_7_6 <= _GEN_8093; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_6 <= 1'h0;
      end else begin
        mask_13_7_6 <= _GEN_2029;
      end
    end else begin
      mask_13_7_6 <= _GEN_2029;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_13_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_13_7_7 <= _GEN_12253;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_13_7_7 <= _GEN_8157; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hd == line_mask_clean_line_1) begin
        mask_13_7_7 <= 1'h0;
      end else begin
        mask_13_7_7 <= _GEN_2045;
      end
    end else begin
      mask_13_7_7 <= _GEN_2045;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_14_0_0 <= _GEN_8222;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_14_0_0 <= _GEN_4126; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_0 <= 1'h0;
      end else begin
        mask_14_0_0 <= _GEN_1038;
      end
    end else begin
      mask_14_0_0 <= _GEN_1038;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_14_0_1 <= _GEN_8286;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_14_0_1 <= _GEN_4190; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_1 <= 1'h0;
      end else begin
        mask_14_0_1 <= _GEN_1054;
      end
    end else begin
      mask_14_0_1 <= _GEN_1054;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_14_0_2 <= _GEN_8350;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_14_0_2 <= _GEN_4254; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_2 <= 1'h0;
      end else begin
        mask_14_0_2 <= _GEN_1070;
      end
    end else begin
      mask_14_0_2 <= _GEN_1070;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_14_0_3 <= _GEN_8414;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_14_0_3 <= _GEN_4318; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_3 <= 1'h0;
      end else begin
        mask_14_0_3 <= _GEN_1086;
      end
    end else begin
      mask_14_0_3 <= _GEN_1086;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_14_0_4 <= _GEN_8478;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_14_0_4 <= _GEN_4382; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_4 <= 1'h0;
      end else begin
        mask_14_0_4 <= _GEN_1102;
      end
    end else begin
      mask_14_0_4 <= _GEN_1102;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_14_0_5 <= _GEN_8542;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_14_0_5 <= _GEN_4446; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_5 <= 1'h0;
      end else begin
        mask_14_0_5 <= _GEN_1118;
      end
    end else begin
      mask_14_0_5 <= _GEN_1118;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_14_0_6 <= _GEN_8606;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_14_0_6 <= _GEN_4510; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_6 <= 1'h0;
      end else begin
        mask_14_0_6 <= _GEN_1134;
      end
    end else begin
      mask_14_0_6 <= _GEN_1134;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_14_0_7 <= _GEN_8670;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_14_0_7 <= _GEN_4574; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_0_7 <= 1'h0;
      end else begin
        mask_14_0_7 <= _GEN_1150;
      end
    end else begin
      mask_14_0_7 <= _GEN_1150;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_14_1_0 <= _GEN_8734;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_14_1_0 <= _GEN_4638; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_0 <= 1'h0;
      end else begin
        mask_14_1_0 <= _GEN_1166;
      end
    end else begin
      mask_14_1_0 <= _GEN_1166;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_14_1_1 <= _GEN_8798;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_14_1_1 <= _GEN_4702; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_1 <= 1'h0;
      end else begin
        mask_14_1_1 <= _GEN_1182;
      end
    end else begin
      mask_14_1_1 <= _GEN_1182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_14_1_2 <= _GEN_8862;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_14_1_2 <= _GEN_4766; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_2 <= 1'h0;
      end else begin
        mask_14_1_2 <= _GEN_1198;
      end
    end else begin
      mask_14_1_2 <= _GEN_1198;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_14_1_3 <= _GEN_8926;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_14_1_3 <= _GEN_4830; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_3 <= 1'h0;
      end else begin
        mask_14_1_3 <= _GEN_1214;
      end
    end else begin
      mask_14_1_3 <= _GEN_1214;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_14_1_4 <= _GEN_8990;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_14_1_4 <= _GEN_4894; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_4 <= 1'h0;
      end else begin
        mask_14_1_4 <= _GEN_1230;
      end
    end else begin
      mask_14_1_4 <= _GEN_1230;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_14_1_5 <= _GEN_9054;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_14_1_5 <= _GEN_4958; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_5 <= 1'h0;
      end else begin
        mask_14_1_5 <= _GEN_1246;
      end
    end else begin
      mask_14_1_5 <= _GEN_1246;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_14_1_6 <= _GEN_9118;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_14_1_6 <= _GEN_5022; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_6 <= 1'h0;
      end else begin
        mask_14_1_6 <= _GEN_1262;
      end
    end else begin
      mask_14_1_6 <= _GEN_1262;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_14_1_7 <= _GEN_9182;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_14_1_7 <= _GEN_5086; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_1_7 <= 1'h0;
      end else begin
        mask_14_1_7 <= _GEN_1278;
      end
    end else begin
      mask_14_1_7 <= _GEN_1278;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_14_2_0 <= _GEN_9246;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_14_2_0 <= _GEN_5150; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_0 <= 1'h0;
      end else begin
        mask_14_2_0 <= _GEN_1294;
      end
    end else begin
      mask_14_2_0 <= _GEN_1294;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_14_2_1 <= _GEN_9310;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_14_2_1 <= _GEN_5214; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_1 <= 1'h0;
      end else begin
        mask_14_2_1 <= _GEN_1310;
      end
    end else begin
      mask_14_2_1 <= _GEN_1310;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_14_2_2 <= _GEN_9374;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_14_2_2 <= _GEN_5278; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_2 <= 1'h0;
      end else begin
        mask_14_2_2 <= _GEN_1326;
      end
    end else begin
      mask_14_2_2 <= _GEN_1326;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_14_2_3 <= _GEN_9438;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_14_2_3 <= _GEN_5342; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_3 <= 1'h0;
      end else begin
        mask_14_2_3 <= _GEN_1342;
      end
    end else begin
      mask_14_2_3 <= _GEN_1342;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_14_2_4 <= _GEN_9502;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_14_2_4 <= _GEN_5406; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_4 <= 1'h0;
      end else begin
        mask_14_2_4 <= _GEN_1358;
      end
    end else begin
      mask_14_2_4 <= _GEN_1358;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_14_2_5 <= _GEN_9566;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_14_2_5 <= _GEN_5470; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_5 <= 1'h0;
      end else begin
        mask_14_2_5 <= _GEN_1374;
      end
    end else begin
      mask_14_2_5 <= _GEN_1374;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_14_2_6 <= _GEN_9630;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_14_2_6 <= _GEN_5534; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_6 <= 1'h0;
      end else begin
        mask_14_2_6 <= _GEN_1390;
      end
    end else begin
      mask_14_2_6 <= _GEN_1390;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_14_2_7 <= _GEN_9694;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_14_2_7 <= _GEN_5598; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_2_7 <= 1'h0;
      end else begin
        mask_14_2_7 <= _GEN_1406;
      end
    end else begin
      mask_14_2_7 <= _GEN_1406;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_14_3_0 <= _GEN_9758;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_14_3_0 <= _GEN_5662; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_0 <= 1'h0;
      end else begin
        mask_14_3_0 <= _GEN_1422;
      end
    end else begin
      mask_14_3_0 <= _GEN_1422;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_14_3_1 <= _GEN_9822;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_14_3_1 <= _GEN_5726; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_1 <= 1'h0;
      end else begin
        mask_14_3_1 <= _GEN_1438;
      end
    end else begin
      mask_14_3_1 <= _GEN_1438;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_14_3_2 <= _GEN_9886;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_14_3_2 <= _GEN_5790; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_2 <= 1'h0;
      end else begin
        mask_14_3_2 <= _GEN_1454;
      end
    end else begin
      mask_14_3_2 <= _GEN_1454;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_14_3_3 <= _GEN_9950;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_14_3_3 <= _GEN_5854; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_3 <= 1'h0;
      end else begin
        mask_14_3_3 <= _GEN_1470;
      end
    end else begin
      mask_14_3_3 <= _GEN_1470;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_14_3_4 <= _GEN_10014;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_14_3_4 <= _GEN_5918; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_4 <= 1'h0;
      end else begin
        mask_14_3_4 <= _GEN_1486;
      end
    end else begin
      mask_14_3_4 <= _GEN_1486;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_14_3_5 <= _GEN_10078;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_14_3_5 <= _GEN_5982; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_5 <= 1'h0;
      end else begin
        mask_14_3_5 <= _GEN_1502;
      end
    end else begin
      mask_14_3_5 <= _GEN_1502;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_14_3_6 <= _GEN_10142;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_14_3_6 <= _GEN_6046; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_6 <= 1'h0;
      end else begin
        mask_14_3_6 <= _GEN_1518;
      end
    end else begin
      mask_14_3_6 <= _GEN_1518;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_14_3_7 <= _GEN_10206;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_14_3_7 <= _GEN_6110; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_3_7 <= 1'h0;
      end else begin
        mask_14_3_7 <= _GEN_1534;
      end
    end else begin
      mask_14_3_7 <= _GEN_1534;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_14_4_0 <= _GEN_10270;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_14_4_0 <= _GEN_6174; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_0 <= 1'h0;
      end else begin
        mask_14_4_0 <= _GEN_1550;
      end
    end else begin
      mask_14_4_0 <= _GEN_1550;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_14_4_1 <= _GEN_10334;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_14_4_1 <= _GEN_6238; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_1 <= 1'h0;
      end else begin
        mask_14_4_1 <= _GEN_1566;
      end
    end else begin
      mask_14_4_1 <= _GEN_1566;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_14_4_2 <= _GEN_10398;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_14_4_2 <= _GEN_6302; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_2 <= 1'h0;
      end else begin
        mask_14_4_2 <= _GEN_1582;
      end
    end else begin
      mask_14_4_2 <= _GEN_1582;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_14_4_3 <= _GEN_10462;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_14_4_3 <= _GEN_6366; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_3 <= 1'h0;
      end else begin
        mask_14_4_3 <= _GEN_1598;
      end
    end else begin
      mask_14_4_3 <= _GEN_1598;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_14_4_4 <= _GEN_10526;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_14_4_4 <= _GEN_6430; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_4 <= 1'h0;
      end else begin
        mask_14_4_4 <= _GEN_1614;
      end
    end else begin
      mask_14_4_4 <= _GEN_1614;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_14_4_5 <= _GEN_10590;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_14_4_5 <= _GEN_6494; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_5 <= 1'h0;
      end else begin
        mask_14_4_5 <= _GEN_1630;
      end
    end else begin
      mask_14_4_5 <= _GEN_1630;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_14_4_6 <= _GEN_10654;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_14_4_6 <= _GEN_6558; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_6 <= 1'h0;
      end else begin
        mask_14_4_6 <= _GEN_1646;
      end
    end else begin
      mask_14_4_6 <= _GEN_1646;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_14_4_7 <= _GEN_10718;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_14_4_7 <= _GEN_6622; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_4_7 <= 1'h0;
      end else begin
        mask_14_4_7 <= _GEN_1662;
      end
    end else begin
      mask_14_4_7 <= _GEN_1662;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_14_5_0 <= _GEN_10782;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_14_5_0 <= _GEN_6686; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_0 <= 1'h0;
      end else begin
        mask_14_5_0 <= _GEN_1678;
      end
    end else begin
      mask_14_5_0 <= _GEN_1678;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_14_5_1 <= _GEN_10846;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_14_5_1 <= _GEN_6750; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_1 <= 1'h0;
      end else begin
        mask_14_5_1 <= _GEN_1694;
      end
    end else begin
      mask_14_5_1 <= _GEN_1694;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_14_5_2 <= _GEN_10910;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_14_5_2 <= _GEN_6814; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_2 <= 1'h0;
      end else begin
        mask_14_5_2 <= _GEN_1710;
      end
    end else begin
      mask_14_5_2 <= _GEN_1710;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_14_5_3 <= _GEN_10974;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_14_5_3 <= _GEN_6878; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_3 <= 1'h0;
      end else begin
        mask_14_5_3 <= _GEN_1726;
      end
    end else begin
      mask_14_5_3 <= _GEN_1726;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_14_5_4 <= _GEN_11038;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_14_5_4 <= _GEN_6942; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_4 <= 1'h0;
      end else begin
        mask_14_5_4 <= _GEN_1742;
      end
    end else begin
      mask_14_5_4 <= _GEN_1742;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_14_5_5 <= _GEN_11102;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_14_5_5 <= _GEN_7006; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_5 <= 1'h0;
      end else begin
        mask_14_5_5 <= _GEN_1758;
      end
    end else begin
      mask_14_5_5 <= _GEN_1758;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_14_5_6 <= _GEN_11166;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_14_5_6 <= _GEN_7070; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_6 <= 1'h0;
      end else begin
        mask_14_5_6 <= _GEN_1774;
      end
    end else begin
      mask_14_5_6 <= _GEN_1774;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_14_5_7 <= _GEN_11230;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_14_5_7 <= _GEN_7134; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_5_7 <= 1'h0;
      end else begin
        mask_14_5_7 <= _GEN_1790;
      end
    end else begin
      mask_14_5_7 <= _GEN_1790;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_14_6_0 <= _GEN_11294;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_14_6_0 <= _GEN_7198; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_0 <= 1'h0;
      end else begin
        mask_14_6_0 <= _GEN_1806;
      end
    end else begin
      mask_14_6_0 <= _GEN_1806;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_14_6_1 <= _GEN_11358;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_14_6_1 <= _GEN_7262; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_1 <= 1'h0;
      end else begin
        mask_14_6_1 <= _GEN_1822;
      end
    end else begin
      mask_14_6_1 <= _GEN_1822;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_14_6_2 <= _GEN_11422;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_14_6_2 <= _GEN_7326; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_2 <= 1'h0;
      end else begin
        mask_14_6_2 <= _GEN_1838;
      end
    end else begin
      mask_14_6_2 <= _GEN_1838;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_14_6_3 <= _GEN_11486;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_14_6_3 <= _GEN_7390; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_3 <= 1'h0;
      end else begin
        mask_14_6_3 <= _GEN_1854;
      end
    end else begin
      mask_14_6_3 <= _GEN_1854;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_14_6_4 <= _GEN_11550;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_14_6_4 <= _GEN_7454; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_4 <= 1'h0;
      end else begin
        mask_14_6_4 <= _GEN_1870;
      end
    end else begin
      mask_14_6_4 <= _GEN_1870;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_14_6_5 <= _GEN_11614;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_14_6_5 <= _GEN_7518; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_5 <= 1'h0;
      end else begin
        mask_14_6_5 <= _GEN_1886;
      end
    end else begin
      mask_14_6_5 <= _GEN_1886;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_14_6_6 <= _GEN_11678;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_14_6_6 <= _GEN_7582; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_6 <= 1'h0;
      end else begin
        mask_14_6_6 <= _GEN_1902;
      end
    end else begin
      mask_14_6_6 <= _GEN_1902;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_14_6_7 <= _GEN_11742;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_14_6_7 <= _GEN_7646; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_6_7 <= 1'h0;
      end else begin
        mask_14_6_7 <= _GEN_1918;
      end
    end else begin
      mask_14_6_7 <= _GEN_1918;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_14_7_0 <= _GEN_11806;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_14_7_0 <= _GEN_7710; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_0 <= 1'h0;
      end else begin
        mask_14_7_0 <= _GEN_1934;
      end
    end else begin
      mask_14_7_0 <= _GEN_1934;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_14_7_1 <= _GEN_11870;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_14_7_1 <= _GEN_7774; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_1 <= 1'h0;
      end else begin
        mask_14_7_1 <= _GEN_1950;
      end
    end else begin
      mask_14_7_1 <= _GEN_1950;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_14_7_2 <= _GEN_11934;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_14_7_2 <= _GEN_7838; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_2 <= 1'h0;
      end else begin
        mask_14_7_2 <= _GEN_1966;
      end
    end else begin
      mask_14_7_2 <= _GEN_1966;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_14_7_3 <= _GEN_11998;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_14_7_3 <= _GEN_7902; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_3 <= 1'h0;
      end else begin
        mask_14_7_3 <= _GEN_1982;
      end
    end else begin
      mask_14_7_3 <= _GEN_1982;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_14_7_4 <= _GEN_12062;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_14_7_4 <= _GEN_7966; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_4 <= 1'h0;
      end else begin
        mask_14_7_4 <= _GEN_1998;
      end
    end else begin
      mask_14_7_4 <= _GEN_1998;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_14_7_5 <= _GEN_12126;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_14_7_5 <= _GEN_8030; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_5 <= 1'h0;
      end else begin
        mask_14_7_5 <= _GEN_2014;
      end
    end else begin
      mask_14_7_5 <= _GEN_2014;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_14_7_6 <= _GEN_12190;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_14_7_6 <= _GEN_8094; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_6 <= 1'h0;
      end else begin
        mask_14_7_6 <= _GEN_2030;
      end
    end else begin
      mask_14_7_6 <= _GEN_2030;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_14_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_14_7_7 <= _GEN_12254;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_14_7_7 <= _GEN_8158; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'he == line_mask_clean_line_1) begin
        mask_14_7_7 <= 1'h0;
      end else begin
        mask_14_7_7 <= _GEN_2046;
      end
    end else begin
      mask_14_7_7 <= _GEN_2046;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_0 <= 1'h0;
    end else if (wen_64) begin // @[Sbuffer.scala 160:18]
      mask_15_0_0 <= _GEN_8223;
    end else if (wen) begin // @[Sbuffer.scala 134:17]
      mask_15_0_0 <= _GEN_4127; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_0 <= 1'h0;
      end else begin
        mask_15_0_0 <= _GEN_1039;
      end
    end else begin
      mask_15_0_0 <= _GEN_1039;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_1 <= 1'h0;
    end else if (wen_65) begin // @[Sbuffer.scala 160:18]
      mask_15_0_1 <= _GEN_8287;
    end else if (wen_1) begin // @[Sbuffer.scala 134:17]
      mask_15_0_1 <= _GEN_4191; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_1 <= 1'h0;
      end else begin
        mask_15_0_1 <= _GEN_1055;
      end
    end else begin
      mask_15_0_1 <= _GEN_1055;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_2 <= 1'h0;
    end else if (wen_66) begin // @[Sbuffer.scala 160:18]
      mask_15_0_2 <= _GEN_8351;
    end else if (wen_2) begin // @[Sbuffer.scala 134:17]
      mask_15_0_2 <= _GEN_4255; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_2 <= 1'h0;
      end else begin
        mask_15_0_2 <= _GEN_1071;
      end
    end else begin
      mask_15_0_2 <= _GEN_1071;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_3 <= 1'h0;
    end else if (wen_67) begin // @[Sbuffer.scala 160:18]
      mask_15_0_3 <= _GEN_8415;
    end else if (wen_3) begin // @[Sbuffer.scala 134:17]
      mask_15_0_3 <= _GEN_4319; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_3 <= 1'h0;
      end else begin
        mask_15_0_3 <= _GEN_1087;
      end
    end else begin
      mask_15_0_3 <= _GEN_1087;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_4 <= 1'h0;
    end else if (wen_68) begin // @[Sbuffer.scala 160:18]
      mask_15_0_4 <= _GEN_8479;
    end else if (wen_4) begin // @[Sbuffer.scala 134:17]
      mask_15_0_4 <= _GEN_4383; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_4 <= 1'h0;
      end else begin
        mask_15_0_4 <= _GEN_1103;
      end
    end else begin
      mask_15_0_4 <= _GEN_1103;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_5 <= 1'h0;
    end else if (wen_69) begin // @[Sbuffer.scala 160:18]
      mask_15_0_5 <= _GEN_8543;
    end else if (wen_5) begin // @[Sbuffer.scala 134:17]
      mask_15_0_5 <= _GEN_4447; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_5 <= 1'h0;
      end else begin
        mask_15_0_5 <= _GEN_1119;
      end
    end else begin
      mask_15_0_5 <= _GEN_1119;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_6 <= 1'h0;
    end else if (wen_70) begin // @[Sbuffer.scala 160:18]
      mask_15_0_6 <= _GEN_8607;
    end else if (wen_6) begin // @[Sbuffer.scala 134:17]
      mask_15_0_6 <= _GEN_4511; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_6 <= 1'h0;
      end else begin
        mask_15_0_6 <= _GEN_1135;
      end
    end else begin
      mask_15_0_6 <= _GEN_1135;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_0_7 <= 1'h0;
    end else if (wen_71) begin // @[Sbuffer.scala 160:18]
      mask_15_0_7 <= _GEN_8671;
    end else if (wen_7) begin // @[Sbuffer.scala 134:17]
      mask_15_0_7 <= _GEN_4575; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_0_7 <= 1'h0;
      end else begin
        mask_15_0_7 <= _GEN_1151;
      end
    end else begin
      mask_15_0_7 <= _GEN_1151;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_0 <= 1'h0;
    end else if (wen_72) begin // @[Sbuffer.scala 160:18]
      mask_15_1_0 <= _GEN_8735;
    end else if (wen_8) begin // @[Sbuffer.scala 134:17]
      mask_15_1_0 <= _GEN_4639; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_0 <= 1'h0;
      end else begin
        mask_15_1_0 <= _GEN_1167;
      end
    end else begin
      mask_15_1_0 <= _GEN_1167;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_1 <= 1'h0;
    end else if (wen_73) begin // @[Sbuffer.scala 160:18]
      mask_15_1_1 <= _GEN_8799;
    end else if (wen_9) begin // @[Sbuffer.scala 134:17]
      mask_15_1_1 <= _GEN_4703; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_1 <= 1'h0;
      end else begin
        mask_15_1_1 <= _GEN_1183;
      end
    end else begin
      mask_15_1_1 <= _GEN_1183;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_2 <= 1'h0;
    end else if (wen_74) begin // @[Sbuffer.scala 160:18]
      mask_15_1_2 <= _GEN_8863;
    end else if (wen_10) begin // @[Sbuffer.scala 134:17]
      mask_15_1_2 <= _GEN_4767; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_2 <= 1'h0;
      end else begin
        mask_15_1_2 <= _GEN_1199;
      end
    end else begin
      mask_15_1_2 <= _GEN_1199;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_3 <= 1'h0;
    end else if (wen_75) begin // @[Sbuffer.scala 160:18]
      mask_15_1_3 <= _GEN_8927;
    end else if (wen_11) begin // @[Sbuffer.scala 134:17]
      mask_15_1_3 <= _GEN_4831; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_3 <= 1'h0;
      end else begin
        mask_15_1_3 <= _GEN_1215;
      end
    end else begin
      mask_15_1_3 <= _GEN_1215;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_4 <= 1'h0;
    end else if (wen_76) begin // @[Sbuffer.scala 160:18]
      mask_15_1_4 <= _GEN_8991;
    end else if (wen_12) begin // @[Sbuffer.scala 134:17]
      mask_15_1_4 <= _GEN_4895; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_4 <= 1'h0;
      end else begin
        mask_15_1_4 <= _GEN_1231;
      end
    end else begin
      mask_15_1_4 <= _GEN_1231;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_5 <= 1'h0;
    end else if (wen_77) begin // @[Sbuffer.scala 160:18]
      mask_15_1_5 <= _GEN_9055;
    end else if (wen_13) begin // @[Sbuffer.scala 134:17]
      mask_15_1_5 <= _GEN_4959; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_5 <= 1'h0;
      end else begin
        mask_15_1_5 <= _GEN_1247;
      end
    end else begin
      mask_15_1_5 <= _GEN_1247;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_6 <= 1'h0;
    end else if (wen_78) begin // @[Sbuffer.scala 160:18]
      mask_15_1_6 <= _GEN_9119;
    end else if (wen_14) begin // @[Sbuffer.scala 134:17]
      mask_15_1_6 <= _GEN_5023; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_6 <= 1'h0;
      end else begin
        mask_15_1_6 <= _GEN_1263;
      end
    end else begin
      mask_15_1_6 <= _GEN_1263;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_1_7 <= 1'h0;
    end else if (wen_79) begin // @[Sbuffer.scala 160:18]
      mask_15_1_7 <= _GEN_9183;
    end else if (wen_15) begin // @[Sbuffer.scala 134:17]
      mask_15_1_7 <= _GEN_5087; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_1_7 <= 1'h0;
      end else begin
        mask_15_1_7 <= _GEN_1279;
      end
    end else begin
      mask_15_1_7 <= _GEN_1279;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_0 <= 1'h0;
    end else if (wen_80) begin // @[Sbuffer.scala 160:18]
      mask_15_2_0 <= _GEN_9247;
    end else if (wen_16) begin // @[Sbuffer.scala 134:17]
      mask_15_2_0 <= _GEN_5151; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_0 <= 1'h0;
      end else begin
        mask_15_2_0 <= _GEN_1295;
      end
    end else begin
      mask_15_2_0 <= _GEN_1295;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_1 <= 1'h0;
    end else if (wen_81) begin // @[Sbuffer.scala 160:18]
      mask_15_2_1 <= _GEN_9311;
    end else if (wen_17) begin // @[Sbuffer.scala 134:17]
      mask_15_2_1 <= _GEN_5215; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_1 <= 1'h0;
      end else begin
        mask_15_2_1 <= _GEN_1311;
      end
    end else begin
      mask_15_2_1 <= _GEN_1311;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_2 <= 1'h0;
    end else if (wen_82) begin // @[Sbuffer.scala 160:18]
      mask_15_2_2 <= _GEN_9375;
    end else if (wen_18) begin // @[Sbuffer.scala 134:17]
      mask_15_2_2 <= _GEN_5279; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_2 <= 1'h0;
      end else begin
        mask_15_2_2 <= _GEN_1327;
      end
    end else begin
      mask_15_2_2 <= _GEN_1327;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_3 <= 1'h0;
    end else if (wen_83) begin // @[Sbuffer.scala 160:18]
      mask_15_2_3 <= _GEN_9439;
    end else if (wen_19) begin // @[Sbuffer.scala 134:17]
      mask_15_2_3 <= _GEN_5343; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_3 <= 1'h0;
      end else begin
        mask_15_2_3 <= _GEN_1343;
      end
    end else begin
      mask_15_2_3 <= _GEN_1343;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_4 <= 1'h0;
    end else if (wen_84) begin // @[Sbuffer.scala 160:18]
      mask_15_2_4 <= _GEN_9503;
    end else if (wen_20) begin // @[Sbuffer.scala 134:17]
      mask_15_2_4 <= _GEN_5407; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_4 <= 1'h0;
      end else begin
        mask_15_2_4 <= _GEN_1359;
      end
    end else begin
      mask_15_2_4 <= _GEN_1359;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_5 <= 1'h0;
    end else if (wen_85) begin // @[Sbuffer.scala 160:18]
      mask_15_2_5 <= _GEN_9567;
    end else if (wen_21) begin // @[Sbuffer.scala 134:17]
      mask_15_2_5 <= _GEN_5471; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_5 <= 1'h0;
      end else begin
        mask_15_2_5 <= _GEN_1375;
      end
    end else begin
      mask_15_2_5 <= _GEN_1375;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_6 <= 1'h0;
    end else if (wen_86) begin // @[Sbuffer.scala 160:18]
      mask_15_2_6 <= _GEN_9631;
    end else if (wen_22) begin // @[Sbuffer.scala 134:17]
      mask_15_2_6 <= _GEN_5535; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_6 <= 1'h0;
      end else begin
        mask_15_2_6 <= _GEN_1391;
      end
    end else begin
      mask_15_2_6 <= _GEN_1391;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_2_7 <= 1'h0;
    end else if (wen_87) begin // @[Sbuffer.scala 160:18]
      mask_15_2_7 <= _GEN_9695;
    end else if (wen_23) begin // @[Sbuffer.scala 134:17]
      mask_15_2_7 <= _GEN_5599; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_2_7 <= 1'h0;
      end else begin
        mask_15_2_7 <= _GEN_1407;
      end
    end else begin
      mask_15_2_7 <= _GEN_1407;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_0 <= 1'h0;
    end else if (wen_88) begin // @[Sbuffer.scala 160:18]
      mask_15_3_0 <= _GEN_9759;
    end else if (wen_24) begin // @[Sbuffer.scala 134:17]
      mask_15_3_0 <= _GEN_5663; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_0 <= 1'h0;
      end else begin
        mask_15_3_0 <= _GEN_1423;
      end
    end else begin
      mask_15_3_0 <= _GEN_1423;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_1 <= 1'h0;
    end else if (wen_89) begin // @[Sbuffer.scala 160:18]
      mask_15_3_1 <= _GEN_9823;
    end else if (wen_25) begin // @[Sbuffer.scala 134:17]
      mask_15_3_1 <= _GEN_5727; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_1 <= 1'h0;
      end else begin
        mask_15_3_1 <= _GEN_1439;
      end
    end else begin
      mask_15_3_1 <= _GEN_1439;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_2 <= 1'h0;
    end else if (wen_90) begin // @[Sbuffer.scala 160:18]
      mask_15_3_2 <= _GEN_9887;
    end else if (wen_26) begin // @[Sbuffer.scala 134:17]
      mask_15_3_2 <= _GEN_5791; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_2 <= 1'h0;
      end else begin
        mask_15_3_2 <= _GEN_1455;
      end
    end else begin
      mask_15_3_2 <= _GEN_1455;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_3 <= 1'h0;
    end else if (wen_91) begin // @[Sbuffer.scala 160:18]
      mask_15_3_3 <= _GEN_9951;
    end else if (wen_27) begin // @[Sbuffer.scala 134:17]
      mask_15_3_3 <= _GEN_5855; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_3 <= 1'h0;
      end else begin
        mask_15_3_3 <= _GEN_1471;
      end
    end else begin
      mask_15_3_3 <= _GEN_1471;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_4 <= 1'h0;
    end else if (wen_92) begin // @[Sbuffer.scala 160:18]
      mask_15_3_4 <= _GEN_10015;
    end else if (wen_28) begin // @[Sbuffer.scala 134:17]
      mask_15_3_4 <= _GEN_5919; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_4 <= 1'h0;
      end else begin
        mask_15_3_4 <= _GEN_1487;
      end
    end else begin
      mask_15_3_4 <= _GEN_1487;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_5 <= 1'h0;
    end else if (wen_93) begin // @[Sbuffer.scala 160:18]
      mask_15_3_5 <= _GEN_10079;
    end else if (wen_29) begin // @[Sbuffer.scala 134:17]
      mask_15_3_5 <= _GEN_5983; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_5 <= 1'h0;
      end else begin
        mask_15_3_5 <= _GEN_1503;
      end
    end else begin
      mask_15_3_5 <= _GEN_1503;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_6 <= 1'h0;
    end else if (wen_94) begin // @[Sbuffer.scala 160:18]
      mask_15_3_6 <= _GEN_10143;
    end else if (wen_30) begin // @[Sbuffer.scala 134:17]
      mask_15_3_6 <= _GEN_6047; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_6 <= 1'h0;
      end else begin
        mask_15_3_6 <= _GEN_1519;
      end
    end else begin
      mask_15_3_6 <= _GEN_1519;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_3_7 <= 1'h0;
    end else if (wen_95) begin // @[Sbuffer.scala 160:18]
      mask_15_3_7 <= _GEN_10207;
    end else if (wen_31) begin // @[Sbuffer.scala 134:17]
      mask_15_3_7 <= _GEN_6111; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_3_7 <= 1'h0;
      end else begin
        mask_15_3_7 <= _GEN_1535;
      end
    end else begin
      mask_15_3_7 <= _GEN_1535;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_0 <= 1'h0;
    end else if (wen_96) begin // @[Sbuffer.scala 160:18]
      mask_15_4_0 <= _GEN_10271;
    end else if (wen_32) begin // @[Sbuffer.scala 134:17]
      mask_15_4_0 <= _GEN_6175; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_0 <= 1'h0;
      end else begin
        mask_15_4_0 <= _GEN_1551;
      end
    end else begin
      mask_15_4_0 <= _GEN_1551;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_1 <= 1'h0;
    end else if (wen_97) begin // @[Sbuffer.scala 160:18]
      mask_15_4_1 <= _GEN_10335;
    end else if (wen_33) begin // @[Sbuffer.scala 134:17]
      mask_15_4_1 <= _GEN_6239; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_1 <= 1'h0;
      end else begin
        mask_15_4_1 <= _GEN_1567;
      end
    end else begin
      mask_15_4_1 <= _GEN_1567;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_2 <= 1'h0;
    end else if (wen_98) begin // @[Sbuffer.scala 160:18]
      mask_15_4_2 <= _GEN_10399;
    end else if (wen_34) begin // @[Sbuffer.scala 134:17]
      mask_15_4_2 <= _GEN_6303; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_2 <= 1'h0;
      end else begin
        mask_15_4_2 <= _GEN_1583;
      end
    end else begin
      mask_15_4_2 <= _GEN_1583;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_3 <= 1'h0;
    end else if (wen_99) begin // @[Sbuffer.scala 160:18]
      mask_15_4_3 <= _GEN_10463;
    end else if (wen_35) begin // @[Sbuffer.scala 134:17]
      mask_15_4_3 <= _GEN_6367; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_3 <= 1'h0;
      end else begin
        mask_15_4_3 <= _GEN_1599;
      end
    end else begin
      mask_15_4_3 <= _GEN_1599;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_4 <= 1'h0;
    end else if (wen_100) begin // @[Sbuffer.scala 160:18]
      mask_15_4_4 <= _GEN_10527;
    end else if (wen_36) begin // @[Sbuffer.scala 134:17]
      mask_15_4_4 <= _GEN_6431; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_4 <= 1'h0;
      end else begin
        mask_15_4_4 <= _GEN_1615;
      end
    end else begin
      mask_15_4_4 <= _GEN_1615;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_5 <= 1'h0;
    end else if (wen_101) begin // @[Sbuffer.scala 160:18]
      mask_15_4_5 <= _GEN_10591;
    end else if (wen_37) begin // @[Sbuffer.scala 134:17]
      mask_15_4_5 <= _GEN_6495; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_5 <= 1'h0;
      end else begin
        mask_15_4_5 <= _GEN_1631;
      end
    end else begin
      mask_15_4_5 <= _GEN_1631;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_6 <= 1'h0;
    end else if (wen_102) begin // @[Sbuffer.scala 160:18]
      mask_15_4_6 <= _GEN_10655;
    end else if (wen_38) begin // @[Sbuffer.scala 134:17]
      mask_15_4_6 <= _GEN_6559; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_6 <= 1'h0;
      end else begin
        mask_15_4_6 <= _GEN_1647;
      end
    end else begin
      mask_15_4_6 <= _GEN_1647;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_4_7 <= 1'h0;
    end else if (wen_103) begin // @[Sbuffer.scala 160:18]
      mask_15_4_7 <= _GEN_10719;
    end else if (wen_39) begin // @[Sbuffer.scala 134:17]
      mask_15_4_7 <= _GEN_6623; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_4_7 <= 1'h0;
      end else begin
        mask_15_4_7 <= _GEN_1663;
      end
    end else begin
      mask_15_4_7 <= _GEN_1663;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_0 <= 1'h0;
    end else if (wen_104) begin // @[Sbuffer.scala 160:18]
      mask_15_5_0 <= _GEN_10783;
    end else if (wen_40) begin // @[Sbuffer.scala 134:17]
      mask_15_5_0 <= _GEN_6687; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_0 <= 1'h0;
      end else begin
        mask_15_5_0 <= _GEN_1679;
      end
    end else begin
      mask_15_5_0 <= _GEN_1679;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_1 <= 1'h0;
    end else if (wen_105) begin // @[Sbuffer.scala 160:18]
      mask_15_5_1 <= _GEN_10847;
    end else if (wen_41) begin // @[Sbuffer.scala 134:17]
      mask_15_5_1 <= _GEN_6751; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_1 <= 1'h0;
      end else begin
        mask_15_5_1 <= _GEN_1695;
      end
    end else begin
      mask_15_5_1 <= _GEN_1695;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_2 <= 1'h0;
    end else if (wen_106) begin // @[Sbuffer.scala 160:18]
      mask_15_5_2 <= _GEN_10911;
    end else if (wen_42) begin // @[Sbuffer.scala 134:17]
      mask_15_5_2 <= _GEN_6815; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_2 <= 1'h0;
      end else begin
        mask_15_5_2 <= _GEN_1711;
      end
    end else begin
      mask_15_5_2 <= _GEN_1711;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_3 <= 1'h0;
    end else if (wen_107) begin // @[Sbuffer.scala 160:18]
      mask_15_5_3 <= _GEN_10975;
    end else if (wen_43) begin // @[Sbuffer.scala 134:17]
      mask_15_5_3 <= _GEN_6879; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_3 <= 1'h0;
      end else begin
        mask_15_5_3 <= _GEN_1727;
      end
    end else begin
      mask_15_5_3 <= _GEN_1727;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_4 <= 1'h0;
    end else if (wen_108) begin // @[Sbuffer.scala 160:18]
      mask_15_5_4 <= _GEN_11039;
    end else if (wen_44) begin // @[Sbuffer.scala 134:17]
      mask_15_5_4 <= _GEN_6943; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_4 <= 1'h0;
      end else begin
        mask_15_5_4 <= _GEN_1743;
      end
    end else begin
      mask_15_5_4 <= _GEN_1743;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_5 <= 1'h0;
    end else if (wen_109) begin // @[Sbuffer.scala 160:18]
      mask_15_5_5 <= _GEN_11103;
    end else if (wen_45) begin // @[Sbuffer.scala 134:17]
      mask_15_5_5 <= _GEN_7007; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_5 <= 1'h0;
      end else begin
        mask_15_5_5 <= _GEN_1759;
      end
    end else begin
      mask_15_5_5 <= _GEN_1759;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_6 <= 1'h0;
    end else if (wen_110) begin // @[Sbuffer.scala 160:18]
      mask_15_5_6 <= _GEN_11167;
    end else if (wen_46) begin // @[Sbuffer.scala 134:17]
      mask_15_5_6 <= _GEN_7071; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_6 <= 1'h0;
      end else begin
        mask_15_5_6 <= _GEN_1775;
      end
    end else begin
      mask_15_5_6 <= _GEN_1775;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_5_7 <= 1'h0;
    end else if (wen_111) begin // @[Sbuffer.scala 160:18]
      mask_15_5_7 <= _GEN_11231;
    end else if (wen_47) begin // @[Sbuffer.scala 134:17]
      mask_15_5_7 <= _GEN_7135; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_5_7 <= 1'h0;
      end else begin
        mask_15_5_7 <= _GEN_1791;
      end
    end else begin
      mask_15_5_7 <= _GEN_1791;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_0 <= 1'h0;
    end else if (wen_112) begin // @[Sbuffer.scala 160:18]
      mask_15_6_0 <= _GEN_11295;
    end else if (wen_48) begin // @[Sbuffer.scala 134:17]
      mask_15_6_0 <= _GEN_7199; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_0 <= 1'h0;
      end else begin
        mask_15_6_0 <= _GEN_1807;
      end
    end else begin
      mask_15_6_0 <= _GEN_1807;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_1 <= 1'h0;
    end else if (wen_113) begin // @[Sbuffer.scala 160:18]
      mask_15_6_1 <= _GEN_11359;
    end else if (wen_49) begin // @[Sbuffer.scala 134:17]
      mask_15_6_1 <= _GEN_7263; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_1 <= 1'h0;
      end else begin
        mask_15_6_1 <= _GEN_1823;
      end
    end else begin
      mask_15_6_1 <= _GEN_1823;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_2 <= 1'h0;
    end else if (wen_114) begin // @[Sbuffer.scala 160:18]
      mask_15_6_2 <= _GEN_11423;
    end else if (wen_50) begin // @[Sbuffer.scala 134:17]
      mask_15_6_2 <= _GEN_7327; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_2 <= 1'h0;
      end else begin
        mask_15_6_2 <= _GEN_1839;
      end
    end else begin
      mask_15_6_2 <= _GEN_1839;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_3 <= 1'h0;
    end else if (wen_115) begin // @[Sbuffer.scala 160:18]
      mask_15_6_3 <= _GEN_11487;
    end else if (wen_51) begin // @[Sbuffer.scala 134:17]
      mask_15_6_3 <= _GEN_7391; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_3 <= 1'h0;
      end else begin
        mask_15_6_3 <= _GEN_1855;
      end
    end else begin
      mask_15_6_3 <= _GEN_1855;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_4 <= 1'h0;
    end else if (wen_116) begin // @[Sbuffer.scala 160:18]
      mask_15_6_4 <= _GEN_11551;
    end else if (wen_52) begin // @[Sbuffer.scala 134:17]
      mask_15_6_4 <= _GEN_7455; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_4 <= 1'h0;
      end else begin
        mask_15_6_4 <= _GEN_1871;
      end
    end else begin
      mask_15_6_4 <= _GEN_1871;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_5 <= 1'h0;
    end else if (wen_117) begin // @[Sbuffer.scala 160:18]
      mask_15_6_5 <= _GEN_11615;
    end else if (wen_53) begin // @[Sbuffer.scala 134:17]
      mask_15_6_5 <= _GEN_7519; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_5 <= 1'h0;
      end else begin
        mask_15_6_5 <= _GEN_1887;
      end
    end else begin
      mask_15_6_5 <= _GEN_1887;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_6 <= 1'h0;
    end else if (wen_118) begin // @[Sbuffer.scala 160:18]
      mask_15_6_6 <= _GEN_11679;
    end else if (wen_54) begin // @[Sbuffer.scala 134:17]
      mask_15_6_6 <= _GEN_7583; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_6 <= 1'h0;
      end else begin
        mask_15_6_6 <= _GEN_1903;
      end
    end else begin
      mask_15_6_6 <= _GEN_1903;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_6_7 <= 1'h0;
    end else if (wen_119) begin // @[Sbuffer.scala 160:18]
      mask_15_6_7 <= _GEN_11743;
    end else if (wen_55) begin // @[Sbuffer.scala 134:17]
      mask_15_6_7 <= _GEN_7647; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_6_7 <= 1'h0;
      end else begin
        mask_15_6_7 <= _GEN_1919;
      end
    end else begin
      mask_15_6_7 <= _GEN_1919;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_0 <= 1'h0;
    end else if (wen_120) begin // @[Sbuffer.scala 160:18]
      mask_15_7_0 <= _GEN_11807;
    end else if (wen_56) begin // @[Sbuffer.scala 134:17]
      mask_15_7_0 <= _GEN_7711; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_0 <= 1'h0;
      end else begin
        mask_15_7_0 <= _GEN_1935;
      end
    end else begin
      mask_15_7_0 <= _GEN_1935;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_1 <= 1'h0;
    end else if (wen_121) begin // @[Sbuffer.scala 160:18]
      mask_15_7_1 <= _GEN_11871;
    end else if (wen_57) begin // @[Sbuffer.scala 134:17]
      mask_15_7_1 <= _GEN_7775; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_1 <= 1'h0;
      end else begin
        mask_15_7_1 <= _GEN_1951;
      end
    end else begin
      mask_15_7_1 <= _GEN_1951;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_2 <= 1'h0;
    end else if (wen_122) begin // @[Sbuffer.scala 160:18]
      mask_15_7_2 <= _GEN_11935;
    end else if (wen_58) begin // @[Sbuffer.scala 134:17]
      mask_15_7_2 <= _GEN_7839; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_2 <= 1'h0;
      end else begin
        mask_15_7_2 <= _GEN_1967;
      end
    end else begin
      mask_15_7_2 <= _GEN_1967;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_3 <= 1'h0;
    end else if (wen_123) begin // @[Sbuffer.scala 160:18]
      mask_15_7_3 <= _GEN_11999;
    end else if (wen_59) begin // @[Sbuffer.scala 134:17]
      mask_15_7_3 <= _GEN_7903; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_3 <= 1'h0;
      end else begin
        mask_15_7_3 <= _GEN_1983;
      end
    end else begin
      mask_15_7_3 <= _GEN_1983;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_4 <= 1'h0;
    end else if (wen_124) begin // @[Sbuffer.scala 160:18]
      mask_15_7_4 <= _GEN_12063;
    end else if (wen_60) begin // @[Sbuffer.scala 134:17]
      mask_15_7_4 <= _GEN_7967; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_4 <= 1'h0;
      end else begin
        mask_15_7_4 <= _GEN_1999;
      end
    end else begin
      mask_15_7_4 <= _GEN_1999;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_5 <= 1'h0;
    end else if (wen_125) begin // @[Sbuffer.scala 160:18]
      mask_15_7_5 <= _GEN_12127;
    end else if (wen_61) begin // @[Sbuffer.scala 134:17]
      mask_15_7_5 <= _GEN_8031; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_5 <= 1'h0;
      end else begin
        mask_15_7_5 <= _GEN_2015;
      end
    end else begin
      mask_15_7_5 <= _GEN_2015;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_6 <= 1'h0;
    end else if (wen_126) begin // @[Sbuffer.scala 160:18]
      mask_15_7_6 <= _GEN_12191;
    end else if (wen_62) begin // @[Sbuffer.scala 134:17]
      mask_15_7_6 <= _GEN_8095; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_6 <= 1'h0;
      end else begin
        mask_15_7_6 <= _GEN_2031;
      end
    end else begin
      mask_15_7_6 <= _GEN_2031;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 160:18]
      mask_15_7_7 <= 1'h0;
    end else if (wen_127) begin // @[Sbuffer.scala 160:18]
      mask_15_7_7 <= _GEN_12255;
    end else if (wen_63) begin // @[Sbuffer.scala 134:17]
      mask_15_7_7 <= _GEN_8159; // @[Sbuffer.scala 137:{34,34}]
    end else if (line_mask_clean_valid_1) begin
      if (4'hf == line_mask_clean_line_1) begin
        mask_15_7_7 <= 1'h0;
      end else begin
        mask_15_7_7 <= _GEN_2047;
      end
    end else begin
      mask_15_7_7 <= _GEN_2047;
    end
  end
endmodule