module ValidPLRUWrapper(
  input        clock,
  input        reset,
  input        io_access_0_valid,
  input  [3:0] io_access_0_bits,
  input        io_access_1_valid,
  input  [3:0] io_access_1_bits,
  input        io_access_2_valid,
  input  [3:0] io_access_2_bits,
  input        io_candidateVec_0,
  input        io_candidateVec_1,
  input        io_candidateVec_2,
  input        io_candidateVec_3,
  input        io_candidateVec_4,
  input        io_candidateVec_5,
  input        io_candidateVec_6,
  input        io_candidateVec_7,
  input        io_candidateVec_8,
  input        io_candidateVec_9,
  input        io_candidateVec_10,
  input        io_candidateVec_11,
  input        io_candidateVec_12,
  input        io_candidateVec_13,
  input        io_candidateVec_14,
  input        io_candidateVec_15,
  output [3:0] io_replaceWay
);
  reg [14:0] state_reg; // @[Replacement.scala 168:62]
  wire  _T_1 = io_access_0_valid | io_access_1_valid | io_access_2_valid; // @[package.scala 72:59]
  wire  state_reg_set_left_older = ~io_access_0_bits[3]; // @[Replacement.scala 196:33]
  wire [6:0] state_reg_left_subtree_state = state_reg[13:7]; // @[package.scala 154:13]
  wire [6:0] state_reg_right_subtree_state = state_reg[6:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_1 = ~io_access_0_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_reg_left_subtree_state_1 = state_reg_left_subtree_state[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_1 = state_reg_left_subtree_state[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_2 = ~io_access_0_bits[1]; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state_2 = state_reg_left_subtree_state_1[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_2 = state_reg_left_subtree_state_1[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_4 = ~io_access_0_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_reg_T_5 = state_reg_set_left_older_2 ? state_reg_left_subtree_state_2 : _state_reg_T_4; // @[Replacement.scala 203:16]
  wire  _state_reg_T_9 = state_reg_set_left_older_2 ? _state_reg_T_4 : state_reg_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_10 = {state_reg_set_left_older_2,_state_reg_T_5,_state_reg_T_9}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_11 = state_reg_set_left_older_1 ? state_reg_left_subtree_state_1 : _state_reg_T_10; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_3 = state_reg_right_subtree_state_1[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_3 = state_reg_right_subtree_state_1[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_16 = state_reg_set_left_older_2 ? state_reg_left_subtree_state_3 : _state_reg_T_4; // @[Replacement.scala 203:16]
  wire  _state_reg_T_20 = state_reg_set_left_older_2 ? _state_reg_T_4 : state_reg_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_21 = {state_reg_set_left_older_2,_state_reg_T_16,_state_reg_T_20}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_22 = state_reg_set_left_older_1 ? _state_reg_T_21 : state_reg_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_23 = {state_reg_set_left_older_1,_state_reg_T_11,_state_reg_T_22}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_24 = state_reg_set_left_older ? state_reg_left_subtree_state : _state_reg_T_23; // @[Replacement.scala 203:16]
  wire [2:0] state_reg_left_subtree_state_4 = state_reg_right_subtree_state[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_4 = state_reg_right_subtree_state[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_left_subtree_state_5 = state_reg_left_subtree_state_4[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_5 = state_reg_left_subtree_state_4[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_30 = state_reg_set_left_older_2 ? state_reg_left_subtree_state_5 : _state_reg_T_4; // @[Replacement.scala 203:16]
  wire  _state_reg_T_34 = state_reg_set_left_older_2 ? _state_reg_T_4 : state_reg_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_35 = {state_reg_set_left_older_2,_state_reg_T_30,_state_reg_T_34}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_36 = state_reg_set_left_older_1 ? state_reg_left_subtree_state_4 : _state_reg_T_35; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_6 = state_reg_right_subtree_state_4[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_6 = state_reg_right_subtree_state_4[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_41 = state_reg_set_left_older_2 ? state_reg_left_subtree_state_6 : _state_reg_T_4; // @[Replacement.scala 203:16]
  wire  _state_reg_T_45 = state_reg_set_left_older_2 ? _state_reg_T_4 : state_reg_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_46 = {state_reg_set_left_older_2,_state_reg_T_41,_state_reg_T_45}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_47 = state_reg_set_left_older_1 ? _state_reg_T_46 : state_reg_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_48 = {state_reg_set_left_older_1,_state_reg_T_36,_state_reg_T_47}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_49 = state_reg_set_left_older ? _state_reg_T_48 : state_reg_right_subtree_state; // @[Replacement.scala 206:16]
  wire [14:0] _state_reg_T_50 = {state_reg_set_left_older,_state_reg_T_24,_state_reg_T_49}; // @[Cat.scala 33:92]
  wire [14:0] _state_reg_T_51 = io_access_0_valid ? _state_reg_T_50 : state_reg; // @[Replacement.scala 22:56]
  wire  state_reg_set_left_older_7 = ~io_access_1_bits[3]; // @[Replacement.scala 196:33]
  wire [6:0] state_reg_left_subtree_state_7 = _state_reg_T_51[13:7]; // @[package.scala 154:13]
  wire [6:0] state_reg_right_subtree_state_7 = _state_reg_T_51[6:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_8 = ~io_access_1_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_reg_left_subtree_state_8 = state_reg_left_subtree_state_7[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_8 = state_reg_left_subtree_state_7[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_9 = ~io_access_1_bits[1]; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state_9 = state_reg_left_subtree_state_8[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_9 = state_reg_left_subtree_state_8[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_56 = ~io_access_1_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_reg_T_57 = state_reg_set_left_older_9 ? state_reg_left_subtree_state_9 : _state_reg_T_56; // @[Replacement.scala 203:16]
  wire  _state_reg_T_61 = state_reg_set_left_older_9 ? _state_reg_T_56 : state_reg_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_62 = {state_reg_set_left_older_9,_state_reg_T_57,_state_reg_T_61}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_63 = state_reg_set_left_older_8 ? state_reg_left_subtree_state_8 : _state_reg_T_62; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_10 = state_reg_right_subtree_state_8[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_10 = state_reg_right_subtree_state_8[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_68 = state_reg_set_left_older_9 ? state_reg_left_subtree_state_10 : _state_reg_T_56; // @[Replacement.scala 203:16]
  wire  _state_reg_T_72 = state_reg_set_left_older_9 ? _state_reg_T_56 : state_reg_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_73 = {state_reg_set_left_older_9,_state_reg_T_68,_state_reg_T_72}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_74 = state_reg_set_left_older_8 ? _state_reg_T_73 : state_reg_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_75 = {state_reg_set_left_older_8,_state_reg_T_63,_state_reg_T_74}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_76 = state_reg_set_left_older_7 ? state_reg_left_subtree_state_7 : _state_reg_T_75; // @[Replacement.scala 203:16]
  wire [2:0] state_reg_left_subtree_state_11 = state_reg_right_subtree_state_7[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_11 = state_reg_right_subtree_state_7[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_left_subtree_state_12 = state_reg_left_subtree_state_11[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_12 = state_reg_left_subtree_state_11[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_82 = state_reg_set_left_older_9 ? state_reg_left_subtree_state_12 : _state_reg_T_56; // @[Replacement.scala 203:16]
  wire  _state_reg_T_86 = state_reg_set_left_older_9 ? _state_reg_T_56 : state_reg_right_subtree_state_12; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_87 = {state_reg_set_left_older_9,_state_reg_T_82,_state_reg_T_86}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_88 = state_reg_set_left_older_8 ? state_reg_left_subtree_state_11 : _state_reg_T_87; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_13 = state_reg_right_subtree_state_11[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_13 = state_reg_right_subtree_state_11[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_93 = state_reg_set_left_older_9 ? state_reg_left_subtree_state_13 : _state_reg_T_56; // @[Replacement.scala 203:16]
  wire  _state_reg_T_97 = state_reg_set_left_older_9 ? _state_reg_T_56 : state_reg_right_subtree_state_13; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_98 = {state_reg_set_left_older_9,_state_reg_T_93,_state_reg_T_97}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_99 = state_reg_set_left_older_8 ? _state_reg_T_98 : state_reg_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_100 = {state_reg_set_left_older_8,_state_reg_T_88,_state_reg_T_99}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_101 = state_reg_set_left_older_7 ? _state_reg_T_100 : state_reg_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [14:0] _state_reg_T_102 = {state_reg_set_left_older_7,_state_reg_T_76,_state_reg_T_101}; // @[Cat.scala 33:92]
  wire [14:0] _state_reg_T_103 = io_access_1_valid ? _state_reg_T_102 : _state_reg_T_51; // @[Replacement.scala 22:56]
  wire  state_reg_set_left_older_14 = ~io_access_2_bits[3]; // @[Replacement.scala 196:33]
  wire [6:0] state_reg_left_subtree_state_14 = _state_reg_T_103[13:7]; // @[package.scala 154:13]
  wire [6:0] state_reg_right_subtree_state_14 = _state_reg_T_103[6:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_15 = ~io_access_2_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_reg_left_subtree_state_15 = state_reg_left_subtree_state_14[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_15 = state_reg_left_subtree_state_14[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_set_left_older_16 = ~io_access_2_bits[1]; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state_16 = state_reg_left_subtree_state_15[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_16 = state_reg_left_subtree_state_15[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_108 = ~io_access_2_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_reg_T_109 = state_reg_set_left_older_16 ? state_reg_left_subtree_state_16 : _state_reg_T_108; // @[Replacement.scala 203:16]
  wire  _state_reg_T_113 = state_reg_set_left_older_16 ? _state_reg_T_108 : state_reg_right_subtree_state_16; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_114 = {state_reg_set_left_older_16,_state_reg_T_109,_state_reg_T_113}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_115 = state_reg_set_left_older_15 ? state_reg_left_subtree_state_15 : _state_reg_T_114; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_17 = state_reg_right_subtree_state_15[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_17 = state_reg_right_subtree_state_15[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_120 = state_reg_set_left_older_16 ? state_reg_left_subtree_state_17 : _state_reg_T_108; // @[Replacement.scala 203:16]
  wire  _state_reg_T_124 = state_reg_set_left_older_16 ? _state_reg_T_108 : state_reg_right_subtree_state_17; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_125 = {state_reg_set_left_older_16,_state_reg_T_120,_state_reg_T_124}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_126 = state_reg_set_left_older_15 ? _state_reg_T_125 : state_reg_right_subtree_state_15; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_127 = {state_reg_set_left_older_15,_state_reg_T_115,_state_reg_T_126}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_128 = state_reg_set_left_older_14 ? state_reg_left_subtree_state_14 : _state_reg_T_127; // @[Replacement.scala 203:16]
  wire [2:0] state_reg_left_subtree_state_18 = state_reg_right_subtree_state_14[5:3]; // @[package.scala 154:13]
  wire [2:0] state_reg_right_subtree_state_18 = state_reg_right_subtree_state_14[2:0]; // @[Replacement.scala 198:38]
  wire  state_reg_left_subtree_state_19 = state_reg_left_subtree_state_18[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_19 = state_reg_left_subtree_state_18[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_134 = state_reg_set_left_older_16 ? state_reg_left_subtree_state_19 : _state_reg_T_108; // @[Replacement.scala 203:16]
  wire  _state_reg_T_138 = state_reg_set_left_older_16 ? _state_reg_T_108 : state_reg_right_subtree_state_19; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_139 = {state_reg_set_left_older_16,_state_reg_T_134,_state_reg_T_138}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_140 = state_reg_set_left_older_15 ? state_reg_left_subtree_state_18 : _state_reg_T_139; // @[Replacement.scala 203:16]
  wire  state_reg_left_subtree_state_20 = state_reg_right_subtree_state_18[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state_20 = state_reg_right_subtree_state_18[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_145 = state_reg_set_left_older_16 ? state_reg_left_subtree_state_20 : _state_reg_T_108; // @[Replacement.scala 203:16]
  wire  _state_reg_T_149 = state_reg_set_left_older_16 ? _state_reg_T_108 : state_reg_right_subtree_state_20; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_150 = {state_reg_set_left_older_16,_state_reg_T_145,_state_reg_T_149}; // @[Cat.scala 33:92]
  wire [2:0] _state_reg_T_151 = state_reg_set_left_older_15 ? _state_reg_T_150 : state_reg_right_subtree_state_18; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_152 = {state_reg_set_left_older_15,_state_reg_T_140,_state_reg_T_151}; // @[Cat.scala 33:92]
  wire [6:0] _state_reg_T_153 = state_reg_set_left_older_14 ? _state_reg_T_152 : state_reg_right_subtree_state_14; // @[Replacement.scala 206:16]
  wire [14:0] _state_reg_T_154 = {state_reg_set_left_older_14,_state_reg_T_128,_state_reg_T_153}; // @[Cat.scala 33:92]
  wire  io_replaceWay_left_subtree_older = state_reg[14]; // @[Replacement.scala 564:38]
  wire  io_replaceWay_left_subtree_older_1 = state_reg_left_subtree_state[6]; // @[Replacement.scala 564:38]
  wire  io_replaceWay_left_subtree_older_2 = state_reg_left_subtree_state_1[2]; // @[Replacement.scala 564:38]
  wire  _io_replaceWay_T_5 = io_candidateVec_15 | io_candidateVec_14; // @[Replacement.scala 598:39]
  wire  _GEN_1 = (io_candidateVec_15 | io_candidateVec_14) & io_candidateVec_15; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_left = io_candidateVec_15 & io_candidateVec_14 ? state_reg_left_subtree_state_2 : _GEN_1; // @[Replacement.scala 595:58 597:13]
  wire  _io_replaceWay_T_13 = io_candidateVec_13 | io_candidateVec_12; // @[Replacement.scala 598:39]
  wire  _GEN_3 = (io_candidateVec_13 | io_candidateVec_12) & io_candidateVec_13; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_right = io_candidateVec_13 & io_candidateVec_12 ? state_reg_right_subtree_state_2 : _GEN_3; // @[Replacement.scala 595:58 597:13]
  wire [1:0] _io_replaceWay_res_T_4 = {1'h0,io_replaceWay_left}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_res_T_5 = io_replaceWay_left_subtree_older_2 ? io_replaceWay_left : io_replaceWay_right; // @[Replacement.scala 579:14]
  wire [1:0] _io_replaceWay_res_T_6 = {io_replaceWay_left_subtree_older_2,_io_replaceWay_res_T_5}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_17 = _io_replaceWay_T_5 | _io_replaceWay_T_13; // @[Replacement.scala 582:33]
  wire  _io_replaceWay_res_T_8 = _io_replaceWay_T_5 ? io_replaceWay_left : io_replaceWay_right; // @[Replacement.scala 585:14]
  wire [1:0] _io_replaceWay_res_T_9 = {_io_replaceWay_T_5,_io_replaceWay_res_T_8}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_5 = _io_replaceWay_T_5 | _io_replaceWay_T_13 ? _io_replaceWay_res_T_9 : _io_replaceWay_res_T_4; // @[Replacement.scala 582:53 584:13 574:25]
  wire [1:0] io_replaceWay_left_1 = _io_replaceWay_T_5 & _io_replaceWay_T_13 ? _io_replaceWay_res_T_6 : _GEN_5; // @[Replacement.scala 576:47 578:13]
  wire  io_replaceWay_left_subtree_older_3 = state_reg_right_subtree_state_1[2]; // @[Replacement.scala 564:38]
  wire  _io_replaceWay_T_23 = io_candidateVec_11 | io_candidateVec_10; // @[Replacement.scala 598:39]
  wire  _GEN_7 = (io_candidateVec_11 | io_candidateVec_10) & io_candidateVec_11; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_left_2 = io_candidateVec_11 & io_candidateVec_10 ? state_reg_left_subtree_state_3 : _GEN_7; // @[Replacement.scala 595:58 597:13]
  wire  _io_replaceWay_T_31 = io_candidateVec_9 | io_candidateVec_8; // @[Replacement.scala 598:39]
  wire  _GEN_9 = (io_candidateVec_9 | io_candidateVec_8) & io_candidateVec_9; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_right_1 = io_candidateVec_9 & io_candidateVec_8 ? state_reg_right_subtree_state_3 : _GEN_9; // @[Replacement.scala 595:58 597:13]
  wire [1:0] _io_replaceWay_res_T_14 = {1'h0,io_replaceWay_left_2}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_res_T_15 = io_replaceWay_left_subtree_older_3 ? io_replaceWay_left_2 : io_replaceWay_right_1; // @[Replacement.scala 579:14]
  wire [1:0] _io_replaceWay_res_T_16 = {io_replaceWay_left_subtree_older_3,_io_replaceWay_res_T_15}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_35 = _io_replaceWay_T_23 | _io_replaceWay_T_31; // @[Replacement.scala 582:33]
  wire  _io_replaceWay_res_T_18 = _io_replaceWay_T_23 ? io_replaceWay_left_2 : io_replaceWay_right_1; // @[Replacement.scala 585:14]
  wire [1:0] _io_replaceWay_res_T_19 = {_io_replaceWay_T_23,_io_replaceWay_res_T_18}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_11 = _io_replaceWay_T_23 | _io_replaceWay_T_31 ? _io_replaceWay_res_T_19 : _io_replaceWay_res_T_14; // @[Replacement.scala 582:53 584:13 574:25]
  wire [1:0] io_replaceWay_right_2 = _io_replaceWay_T_23 & _io_replaceWay_T_31 ? _io_replaceWay_res_T_16 : _GEN_11; // @[Replacement.scala 576:47 578:13]
  wire [2:0] _io_replaceWay_res_T_20 = {1'h0,io_replaceWay_left_1}; // @[Cat.scala 33:92]
  wire [1:0] _io_replaceWay_res_T_21 = io_replaceWay_left_subtree_older_1 ? io_replaceWay_left_1 : io_replaceWay_right_2
    ; // @[Replacement.scala 579:14]
  wire [2:0] _io_replaceWay_res_T_22 = {io_replaceWay_left_subtree_older_1,_io_replaceWay_res_T_21}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_37 = _io_replaceWay_T_5 | _io_replaceWay_T_13 | (_io_replaceWay_T_23 | _io_replaceWay_T_31); // @[Replacement.scala 582:33]
  wire [1:0] _io_replaceWay_res_T_24 = _io_replaceWay_T_17 ? io_replaceWay_left_1 : io_replaceWay_right_2; // @[Replacement.scala 585:14]
  wire [2:0] _io_replaceWay_res_T_25 = {_io_replaceWay_T_17,_io_replaceWay_res_T_24}; // @[Cat.scala 33:92]
  wire [2:0] _GEN_13 = _io_replaceWay_T_5 | _io_replaceWay_T_13 | (_io_replaceWay_T_23 | _io_replaceWay_T_31) ?
    _io_replaceWay_res_T_25 : _io_replaceWay_res_T_20; // @[Replacement.scala 582:53 584:13 574:25]
  wire [2:0] io_replaceWay_left_3 = _io_replaceWay_T_17 & _io_replaceWay_T_35 ? _io_replaceWay_res_T_22 : _GEN_13; // @[Replacement.scala 576:47 578:13]
  wire  io_replaceWay_left_subtree_older_4 = state_reg_right_subtree_state[6]; // @[Replacement.scala 564:38]
  wire  io_replaceWay_left_subtree_older_5 = state_reg_left_subtree_state_4[2]; // @[Replacement.scala 564:38]
  wire  _io_replaceWay_T_43 = io_candidateVec_7 | io_candidateVec_6; // @[Replacement.scala 598:39]
  wire  _GEN_15 = (io_candidateVec_7 | io_candidateVec_6) & io_candidateVec_7; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_left_4 = io_candidateVec_7 & io_candidateVec_6 ? state_reg_left_subtree_state_5 : _GEN_15; // @[Replacement.scala 595:58 597:13]
  wire  _io_replaceWay_T_51 = io_candidateVec_5 | io_candidateVec_4; // @[Replacement.scala 598:39]
  wire  _GEN_17 = (io_candidateVec_5 | io_candidateVec_4) & io_candidateVec_5; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_right_3 = io_candidateVec_5 & io_candidateVec_4 ? state_reg_right_subtree_state_5 : _GEN_17; // @[Replacement.scala 595:58 597:13]
  wire [1:0] _io_replaceWay_res_T_30 = {1'h0,io_replaceWay_left_4}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_res_T_31 = io_replaceWay_left_subtree_older_5 ? io_replaceWay_left_4 : io_replaceWay_right_3; // @[Replacement.scala 579:14]
  wire [1:0] _io_replaceWay_res_T_32 = {io_replaceWay_left_subtree_older_5,_io_replaceWay_res_T_31}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_55 = _io_replaceWay_T_43 | _io_replaceWay_T_51; // @[Replacement.scala 582:33]
  wire  _io_replaceWay_res_T_34 = _io_replaceWay_T_43 ? io_replaceWay_left_4 : io_replaceWay_right_3; // @[Replacement.scala 585:14]
  wire [1:0] _io_replaceWay_res_T_35 = {_io_replaceWay_T_43,_io_replaceWay_res_T_34}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_19 = _io_replaceWay_T_43 | _io_replaceWay_T_51 ? _io_replaceWay_res_T_35 : _io_replaceWay_res_T_30; // @[Replacement.scala 582:53 584:13 574:25]
  wire [1:0] io_replaceWay_left_5 = _io_replaceWay_T_43 & _io_replaceWay_T_51 ? _io_replaceWay_res_T_32 : _GEN_19; // @[Replacement.scala 576:47 578:13]
  wire  io_replaceWay_left_subtree_older_6 = state_reg_right_subtree_state_4[2]; // @[Replacement.scala 564:38]
  wire  _io_replaceWay_T_61 = io_candidateVec_3 | io_candidateVec_2; // @[Replacement.scala 598:39]
  wire  _GEN_21 = (io_candidateVec_3 | io_candidateVec_2) & io_candidateVec_3; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_left_6 = io_candidateVec_3 & io_candidateVec_2 ? state_reg_left_subtree_state_6 : _GEN_21; // @[Replacement.scala 595:58 597:13]
  wire  _io_replaceWay_T_69 = io_candidateVec_1 | io_candidateVec_0; // @[Replacement.scala 598:39]
  wire  _GEN_23 = (io_candidateVec_1 | io_candidateVec_0) & io_candidateVec_1; // @[Replacement.scala 598:64 600:13 594:25]
  wire  io_replaceWay_right_4 = io_candidateVec_1 & io_candidateVec_0 ? state_reg_right_subtree_state_6 : _GEN_23; // @[Replacement.scala 595:58 597:13]
  wire [1:0] _io_replaceWay_res_T_40 = {1'h0,io_replaceWay_left_6}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_res_T_41 = io_replaceWay_left_subtree_older_6 ? io_replaceWay_left_6 : io_replaceWay_right_4; // @[Replacement.scala 579:14]
  wire [1:0] _io_replaceWay_res_T_42 = {io_replaceWay_left_subtree_older_6,_io_replaceWay_res_T_41}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_73 = _io_replaceWay_T_61 | _io_replaceWay_T_69; // @[Replacement.scala 582:33]
  wire  _io_replaceWay_res_T_44 = _io_replaceWay_T_61 ? io_replaceWay_left_6 : io_replaceWay_right_4; // @[Replacement.scala 585:14]
  wire [1:0] _io_replaceWay_res_T_45 = {_io_replaceWay_T_61,_io_replaceWay_res_T_44}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_25 = _io_replaceWay_T_61 | _io_replaceWay_T_69 ? _io_replaceWay_res_T_45 : _io_replaceWay_res_T_40; // @[Replacement.scala 582:53 584:13 574:25]
  wire [1:0] io_replaceWay_right_5 = _io_replaceWay_T_61 & _io_replaceWay_T_69 ? _io_replaceWay_res_T_42 : _GEN_25; // @[Replacement.scala 576:47 578:13]
  wire [2:0] _io_replaceWay_res_T_46 = {1'h0,io_replaceWay_left_5}; // @[Cat.scala 33:92]
  wire [1:0] _io_replaceWay_res_T_47 = io_replaceWay_left_subtree_older_4 ? io_replaceWay_left_5 : io_replaceWay_right_5
    ; // @[Replacement.scala 579:14]
  wire [2:0] _io_replaceWay_res_T_48 = {io_replaceWay_left_subtree_older_4,_io_replaceWay_res_T_47}; // @[Cat.scala 33:92]
  wire  _io_replaceWay_T_75 = _io_replaceWay_T_43 | _io_replaceWay_T_51 | (_io_replaceWay_T_61 | _io_replaceWay_T_69); // @[Replacement.scala 582:33]
  wire [1:0] _io_replaceWay_res_T_50 = _io_replaceWay_T_55 ? io_replaceWay_left_5 : io_replaceWay_right_5; // @[Replacement.scala 585:14]
  wire [2:0] _io_replaceWay_res_T_51 = {_io_replaceWay_T_55,_io_replaceWay_res_T_50}; // @[Cat.scala 33:92]
  wire [2:0] _GEN_27 = _io_replaceWay_T_43 | _io_replaceWay_T_51 | (_io_replaceWay_T_61 | _io_replaceWay_T_69) ?
    _io_replaceWay_res_T_51 : _io_replaceWay_res_T_46; // @[Replacement.scala 582:53 584:13 574:25]
  wire [2:0] io_replaceWay_right_6 = _io_replaceWay_T_55 & _io_replaceWay_T_73 ? _io_replaceWay_res_T_48 : _GEN_27; // @[Replacement.scala 576:47 578:13]
  wire [3:0] _io_replaceWay_res_T_52 = {1'h0,io_replaceWay_left_3}; // @[Cat.scala 33:92]
  wire [2:0] _io_replaceWay_res_T_53 = io_replaceWay_left_subtree_older ? io_replaceWay_left_3 : io_replaceWay_right_6; // @[Replacement.scala 579:14]
  wire [3:0] _io_replaceWay_res_T_54 = {io_replaceWay_left_subtree_older,_io_replaceWay_res_T_53}; // @[Cat.scala 33:92]
  wire [2:0] _io_replaceWay_res_T_56 = _io_replaceWay_T_37 ? io_replaceWay_left_3 : io_replaceWay_right_6; // @[Replacement.scala 585:14]
  wire [3:0] _io_replaceWay_res_T_57 = {_io_replaceWay_T_37,_io_replaceWay_res_T_56}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_29 = _io_replaceWay_T_5 | _io_replaceWay_T_13 | (_io_replaceWay_T_23 | _io_replaceWay_T_31) | (
    _io_replaceWay_T_43 | _io_replaceWay_T_51 | (_io_replaceWay_T_61 | _io_replaceWay_T_69)) ? _io_replaceWay_res_T_57
     : _io_replaceWay_res_T_52; // @[Replacement.scala 582:53 584:13 574:25]
  assign io_replaceWay = _io_replaceWay_T_37 & _io_replaceWay_T_75 ? _io_replaceWay_res_T_54 : _GEN_29; // @[Replacement.scala 576:47 578:13]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 175:40]
      state_reg <= 15'h0; // @[Replacement.scala 22:{56,56,56}]
    end else if (_T_1) begin // @[Replacement.scala 168:62]
      if (io_access_2_valid) begin
        state_reg <= _state_reg_T_154;
      end else if (io_access_1_valid) begin
        state_reg <= _state_reg_T_102;
      end else if (io_access_0_valid) begin
        state_reg <= _state_reg_T_50;
      end
    end
  end
endmodule