module Sbuffer(
  input          clock,
  input          reset,
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [35:0]  io_in_0_bits_addr,
  input  [63:0]  io_in_0_bits_data,
  input  [7:0]   io_in_0_bits_mask,
  input  [38:0]  io_in_0_bits_vaddr,
  input          io_in_0_bits_wline,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [35:0]  io_in_1_bits_addr,
  input  [63:0]  io_in_1_bits_data,
  input  [7:0]   io_in_1_bits_mask,
  input  [38:0]  io_in_1_bits_vaddr,
  input          io_in_1_bits_wline,
  input          io_dcache_req_ready,
  output         io_dcache_req_valid,
  output [38:0]  io_dcache_req_bits_vaddr,
  output [35:0]  io_dcache_req_bits_addr,
  output [511:0] io_dcache_req_bits_data,
  output [63:0]  io_dcache_req_bits_mask,
  output [5:0]   io_dcache_req_bits_id,
  input          io_dcache_main_pipe_hit_resp_valid,
  input  [5:0]   io_dcache_main_pipe_hit_resp_bits_id,
  input          io_dcache_refill_hit_resp_valid,
  input  [5:0]   io_dcache_refill_hit_resp_bits_id,
  input          io_dcache_replay_resp_valid,
  input  [5:0]   io_dcache_replay_resp_bits_id,
  input  [38:0]  io_forward_0_vaddr,
  input  [35:0]  io_forward_0_paddr,
  input          io_forward_0_valid,
  output         io_forward_0_forwardMask_0,
  output         io_forward_0_forwardMask_1,
  output         io_forward_0_forwardMask_2,
  output         io_forward_0_forwardMask_3,
  output         io_forward_0_forwardMask_4,
  output         io_forward_0_forwardMask_5,
  output         io_forward_0_forwardMask_6,
  output         io_forward_0_forwardMask_7,
  output [7:0]   io_forward_0_forwardData_0,
  output [7:0]   io_forward_0_forwardData_1,
  output [7:0]   io_forward_0_forwardData_2,
  output [7:0]   io_forward_0_forwardData_3,
  output [7:0]   io_forward_0_forwardData_4,
  output [7:0]   io_forward_0_forwardData_5,
  output [7:0]   io_forward_0_forwardData_6,
  output [7:0]   io_forward_0_forwardData_7,
  output         io_forward_0_matchInvalid,
  input  [38:0]  io_forward_1_vaddr,
  input  [35:0]  io_forward_1_paddr,
  input          io_forward_1_valid,
  output         io_forward_1_forwardMask_0,
  output         io_forward_1_forwardMask_1,
  output         io_forward_1_forwardMask_2,
  output         io_forward_1_forwardMask_3,
  output         io_forward_1_forwardMask_4,
  output         io_forward_1_forwardMask_5,
  output         io_forward_1_forwardMask_6,
  output         io_forward_1_forwardMask_7,
  output [7:0]   io_forward_1_forwardData_0,
  output [7:0]   io_forward_1_forwardData_1,
  output [7:0]   io_forward_1_forwardData_2,
  output [7:0]   io_forward_1_forwardData_3,
  output [7:0]   io_forward_1_forwardData_4,
  output [7:0]   io_forward_1_forwardData_5,
  output [7:0]   io_forward_1_forwardData_6,
  output [7:0]   io_forward_1_forwardData_7,
  output         io_forward_1_matchInvalid,
  input          io_sqempty,
  input          io_flush_valid,
  output         io_flush_empty,
  input  [3:0]   io_csrCtrl_sbuffer_threshold,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value,
  output [5:0]   io_perf_8_value,
  output [5:0]   io_perf_9_value,
  output [5:0]   io_perf_10_value,
  output [5:0]   io_perf_11_value,
  output [5:0]   io_perf_12_value,
  output [5:0]   io_perf_13_value,
  output [5:0]   io_perf_14_value,
  output [5:0]   io_perf_15_value,
  output [5:0]   io_perf_16_value
);
  wire  dataModule_clock; // @[Sbuffer.scala 270:26]
  wire  dataModule_reset; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_writeReq_0_valid; // @[Sbuffer.scala 270:26]
  wire [15:0] dataModule_io_writeReq_0_bits_wvec; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_writeReq_0_bits_mask; // @[Sbuffer.scala 270:26]
  wire [63:0] dataModule_io_writeReq_0_bits_data; // @[Sbuffer.scala 270:26]
  wire [32:0] dataModule_io_writeReq_0_bits_wordOffset; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_writeReq_0_bits_wline; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_writeReq_1_valid; // @[Sbuffer.scala 270:26]
  wire [15:0] dataModule_io_writeReq_1_bits_wvec; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_writeReq_1_bits_mask; // @[Sbuffer.scala 270:26]
  wire [63:0] dataModule_io_writeReq_1_bits_data; // @[Sbuffer.scala 270:26]
  wire [32:0] dataModule_io_writeReq_1_bits_wordOffset; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_writeReq_1_bits_wline; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskFlushReq_0_valid; // @[Sbuffer.scala 270:26]
  wire [15:0] dataModule_io_maskFlushReq_0_bits_wvec; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskFlushReq_1_valid; // @[Sbuffer.scala 270:26]
  wire [15:0] dataModule_io_maskFlushReq_1_bits_wvec; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_0_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_1_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_2_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_3_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_4_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_5_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_6_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_7_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_8_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_9_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_10_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_11_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_12_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_13_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_14_7_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_0_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_1_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_2_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_3_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_4_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_5_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_6_7; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_0; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_1; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_2; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_3; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_4; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_5; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_6; // @[Sbuffer.scala 270:26]
  wire [7:0] dataModule_io_dataOut_15_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_0_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_1_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_2_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_3_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_4_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_5_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_6_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_7_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_8_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_9_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_10_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_11_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_12_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_13_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_14_7_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_0_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_1_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_2_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_3_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_4_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_5_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_6_7; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_0; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_1; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_2; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_3; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_4; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_5; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_6; // @[Sbuffer.scala 270:26]
  wire  dataModule_io_maskOut_15_7_7; // @[Sbuffer.scala 270:26]
  wire  Sbuffer_PLRU_clock; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_reset; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_access_0_valid; // @[Sbuffer.scala 324:20]
  wire [3:0] Sbuffer_PLRU_io_access_0_bits; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_access_1_valid; // @[Sbuffer.scala 324:20]
  wire [3:0] Sbuffer_PLRU_io_access_1_bits; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_access_2_valid; // @[Sbuffer.scala 324:20]
  wire [3:0] Sbuffer_PLRU_io_access_2_bits; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_0; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_1; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_2; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_3; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_4; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_5; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_6; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_7; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_8; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_9; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_10; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_11; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_12; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_13; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_14; // @[Sbuffer.scala 324:20]
  wire  Sbuffer_PLRU_io_candidateVec_15; // @[Sbuffer.scala 324:20]
  wire [3:0] Sbuffer_PLRU_io_replaceWay; // @[Sbuffer.scala 324:20]
  reg [29:0] ptag_0; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_1; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_2; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_3; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_4; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_5; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_6; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_7; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_8; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_9; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_10; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_11; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_12; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_13; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_14; // @[Sbuffer.scala 274:17]
  reg [29:0] ptag_15; // @[Sbuffer.scala 274:17]
  reg [32:0] vtag_0; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_1; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_2; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_3; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_4; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_5; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_6; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_7; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_8; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_9; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_10; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_11; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_12; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_13; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_14; // @[Sbuffer.scala 275:17]
  reg [32:0] vtag_15; // @[Sbuffer.scala 275:17]
  reg [15:0] waitInflightMask_0; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_1; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_2; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_3; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_4; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_5; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_6; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_7; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_8; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_9; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_10; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_11; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_12; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_13; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_14; // @[Sbuffer.scala 277:29]
  reg [15:0] waitInflightMask_15; // @[Sbuffer.scala 277:29]
  reg  stateVec_0_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_0_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_0_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_0_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_1_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_1_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_1_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_1_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_2_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_2_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_2_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_2_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_3_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_3_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_3_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_3_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_4_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_4_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_4_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_4_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_5_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_5_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_5_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_5_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_6_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_6_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_6_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_6_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_7_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_7_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_7_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_7_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_8_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_8_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_8_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_8_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_9_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_9_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_9_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_9_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_10_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_10_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_10_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_10_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_11_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_11_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_11_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_11_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_12_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_12_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_12_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_12_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_13_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_13_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_13_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_13_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_14_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_14_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_14_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_14_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_15_state_valid; // @[Sbuffer.scala 280:25]
  reg  stateVec_15_state_inflight; // @[Sbuffer.scala 280:25]
  reg  stateVec_15_w_timeout; // @[Sbuffer.scala 280:25]
  reg  stateVec_15_w_sameblock_inflight; // @[Sbuffer.scala 280:25]
  reg [20:0] cohCount_0; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_1; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_2; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_3; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_4; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_5; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_6; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_7; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_8; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_9; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_10; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_11; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_12; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_13; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_14; // @[Sbuffer.scala 281:25]
  reg [20:0] cohCount_15; // @[Sbuffer.scala 281:25]
  reg [4:0] missqReplayCount_0; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_1; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_2; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_3; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_4; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_5; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_6; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_7; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_8; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_9; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_10; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_11; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_12; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_13; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_14; // @[Sbuffer.scala 282:33]
  reg [4:0] missqReplayCount_15; // @[Sbuffer.scala 282:33]
  reg [1:0] sbuffer_state; // @[Sbuffer.scala 295:30]
  wire  _candidateVec_T_1 = stateVec_0_state_valid & ~stateVec_0_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_5 = stateVec_1_state_valid & ~stateVec_1_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_9 = stateVec_2_state_valid & ~stateVec_2_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_13 = stateVec_3_state_valid & ~stateVec_3_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_17 = stateVec_4_state_valid & ~stateVec_4_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_21 = stateVec_5_state_valid & ~stateVec_5_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_25 = stateVec_6_state_valid & ~stateVec_6_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_29 = stateVec_7_state_valid & ~stateVec_7_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_33 = stateVec_8_state_valid & ~stateVec_8_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_37 = stateVec_9_state_valid & ~stateVec_9_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_41 = stateVec_10_state_valid & ~stateVec_10_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_45 = stateVec_11_state_valid & ~stateVec_11_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_49 = stateVec_12_state_valid & ~stateVec_12_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_53 = stateVec_13_state_valid & ~stateVec_13_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_57 = stateVec_14_state_valid & ~stateVec_14_state_inflight; // @[Sbuffer.scala 66:50]
  wire  _candidateVec_T_61 = stateVec_15_state_valid & ~stateVec_15_state_inflight; // @[Sbuffer.scala 66:50]
  wire  cohTimeOutMask_0 = cohCount_0[20] & _candidateVec_T_1; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_1 = cohCount_1[20] & _candidateVec_T_5; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_2 = cohCount_2[20] & _candidateVec_T_9; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_3 = cohCount_3[20] & _candidateVec_T_13; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_4 = cohCount_4[20] & _candidateVec_T_17; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_5 = cohCount_5[20] & _candidateVec_T_21; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_6 = cohCount_6[20] & _candidateVec_T_25; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_7 = cohCount_7[20] & _candidateVec_T_29; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_8 = cohCount_8[20] & _candidateVec_T_33; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_9 = cohCount_9[20] & _candidateVec_T_37; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_10 = cohCount_10[20] & _candidateVec_T_41; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_11 = cohCount_11[20] & _candidateVec_T_45; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_12 = cohCount_12[20] & _candidateVec_T_49; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_13 = cohCount_13[20] & _candidateVec_T_53; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_14 = cohCount_14[20] & _candidateVec_T_57; // @[Sbuffer.scala 341:78]
  wire  cohTimeOutMask_15 = cohCount_15[20] & _candidateVec_T_61; // @[Sbuffer.scala 341:78]
  wire [3:0] d_tail = cohTimeOutMask_14 ? 4'he : 4'hf; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail = cohTimeOutMask_14 | cohTimeOutMask_15; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_1 = cohTimeOutMask_13 ? 4'hd : d_tail; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_1 = cohTimeOutMask_13 | f_tail; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_2 = cohTimeOutMask_12 ? 4'hc : d_tail_1; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_2 = cohTimeOutMask_12 | f_tail_1; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_3 = cohTimeOutMask_11 ? 4'hb : d_tail_2; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_3 = cohTimeOutMask_11 | f_tail_2; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_4 = cohTimeOutMask_10 ? 4'ha : d_tail_3; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_4 = cohTimeOutMask_10 | f_tail_3; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_5 = cohTimeOutMask_9 ? 4'h9 : d_tail_4; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_5 = cohTimeOutMask_9 | f_tail_4; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_6 = cohTimeOutMask_8 ? 4'h8 : d_tail_5; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_6 = cohTimeOutMask_8 | f_tail_5; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_7 = cohTimeOutMask_7 ? 4'h7 : d_tail_6; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_7 = cohTimeOutMask_7 | f_tail_6; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_8 = cohTimeOutMask_6 ? 4'h6 : d_tail_7; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_8 = cohTimeOutMask_6 | f_tail_7; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_9 = cohTimeOutMask_5 ? 4'h5 : d_tail_8; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_9 = cohTimeOutMask_5 | f_tail_8; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_10 = cohTimeOutMask_4 ? 4'h4 : d_tail_9; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_10 = cohTimeOutMask_4 | f_tail_9; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_11 = cohTimeOutMask_3 ? 4'h3 : d_tail_10; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_11 = cohTimeOutMask_3 | f_tail_10; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_12 = cohTimeOutMask_2 ? 4'h2 : d_tail_11; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_12 = cohTimeOutMask_2 | f_tail_11; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_13 = cohTimeOutMask_1 ? 4'h1 : d_tail_12; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_13 = cohTimeOutMask_1 | f_tail_12; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] cohTimeOutIdx = cohTimeOutMask_0 ? 4'h0 : d_tail_13; // @[PriorityMuxDefault.scala 46:13]
  wire  cohHasTimeOut = cohTimeOutMask_0 | f_tail_13; // @[PriorityMuxDefault.scala 46:46]
  wire  missqReplayTimeOutMask_0 = missqReplayCount_0[4] & stateVec_0_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_1 = missqReplayCount_1[4] & stateVec_1_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_2 = missqReplayCount_2[4] & stateVec_2_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_3 = missqReplayCount_3[4] & stateVec_3_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_4 = missqReplayCount_4[4] & stateVec_4_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_5 = missqReplayCount_5[4] & stateVec_5_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_6 = missqReplayCount_6[4] & stateVec_6_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_7 = missqReplayCount_7[4] & stateVec_7_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_8 = missqReplayCount_8[4] & stateVec_8_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_9 = missqReplayCount_9[4] & stateVec_9_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_10 = missqReplayCount_10[4] & stateVec_10_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_11 = missqReplayCount_11[4] & stateVec_11_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_12 = missqReplayCount_12[4] & stateVec_12_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_13 = missqReplayCount_13[4] & stateVec_13_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_14 = missqReplayCount_14[4] & stateVec_14_w_timeout; // @[Sbuffer.scala 344:100]
  wire  missqReplayTimeOutMask_15 = missqReplayCount_15[4] & stateVec_15_w_timeout; // @[Sbuffer.scala 344:100]
  wire [3:0] d_tail_14 = missqReplayTimeOutMask_14 ? 4'he : 4'hf; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_14 = missqReplayTimeOutMask_14 | missqReplayTimeOutMask_15; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_15 = missqReplayTimeOutMask_13 ? 4'hd : d_tail_14; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_15 = missqReplayTimeOutMask_13 | f_tail_14; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_16 = missqReplayTimeOutMask_12 ? 4'hc : d_tail_15; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_16 = missqReplayTimeOutMask_12 | f_tail_15; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_17 = missqReplayTimeOutMask_11 ? 4'hb : d_tail_16; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_17 = missqReplayTimeOutMask_11 | f_tail_16; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_18 = missqReplayTimeOutMask_10 ? 4'ha : d_tail_17; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_18 = missqReplayTimeOutMask_10 | f_tail_17; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_19 = missqReplayTimeOutMask_9 ? 4'h9 : d_tail_18; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_19 = missqReplayTimeOutMask_9 | f_tail_18; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_20 = missqReplayTimeOutMask_8 ? 4'h8 : d_tail_19; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_20 = missqReplayTimeOutMask_8 | f_tail_19; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_21 = missqReplayTimeOutMask_7 ? 4'h7 : d_tail_20; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_21 = missqReplayTimeOutMask_7 | f_tail_20; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_22 = missqReplayTimeOutMask_6 ? 4'h6 : d_tail_21; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_22 = missqReplayTimeOutMask_6 | f_tail_21; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_23 = missqReplayTimeOutMask_5 ? 4'h5 : d_tail_22; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_23 = missqReplayTimeOutMask_5 | f_tail_22; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_24 = missqReplayTimeOutMask_4 ? 4'h4 : d_tail_23; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_24 = missqReplayTimeOutMask_4 | f_tail_23; // @[PriorityMuxDefault.scala 46:46]
  wire [3:0] d_tail_25 = missqReplayTimeOutMask_3 ? 4'h3 : d_tail_24; // @[PriorityMuxDefault.scala 46:13]
  wire  f_tail_25 = missqReplayTimeOutMask_3 | f_tail_24; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_26 = missqReplayTimeOutMask_2 | f_tail_25; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_27 = missqReplayTimeOutMask_1 | f_tail_26; // @[PriorityMuxDefault.scala 46:46]
  wire  missqReplayHasTimeOutGen = missqReplayTimeOutMask_0 | f_tail_27; // @[PriorityMuxDefault.scala 46:46]
  reg  missqReplayHasTimeOut_REG; // @[Sbuffer.scala 346:38]
  reg  missqReplayHasTimeOut_REG_1; // @[Sbuffer.scala 346:76]
  wire  missqReplayHasTimeOut = missqReplayHasTimeOut_REG & ~missqReplayHasTimeOut_REG_1; // @[Sbuffer.scala 346:65]
  reg [3:0] missqReplayTimeOutIdx; // @[Reg.scala 19:16]
  wire [3:0] _drainIdx_T = _candidateVec_T_57 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_1 = _candidateVec_T_53 ? 4'hd : _drainIdx_T; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_2 = _candidateVec_T_49 ? 4'hc : _drainIdx_T_1; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_3 = _candidateVec_T_45 ? 4'hb : _drainIdx_T_2; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_4 = _candidateVec_T_41 ? 4'ha : _drainIdx_T_3; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_5 = _candidateVec_T_37 ? 4'h9 : _drainIdx_T_4; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_6 = _candidateVec_T_33 ? 4'h8 : _drainIdx_T_5; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_7 = _candidateVec_T_29 ? 4'h7 : _drainIdx_T_6; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_8 = _candidateVec_T_25 ? 4'h6 : _drainIdx_T_7; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_9 = _candidateVec_T_21 ? 4'h5 : _drainIdx_T_8; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_10 = _candidateVec_T_17 ? 4'h4 : _drainIdx_T_9; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_11 = _candidateVec_T_13 ? 4'h3 : _drainIdx_T_10; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_12 = _candidateVec_T_9 ? 4'h2 : _drainIdx_T_11; // @[Mux.scala 47:70]
  wire [3:0] _drainIdx_T_13 = _candidateVec_T_5 ? 4'h1 : _drainIdx_T_12; // @[Mux.scala 47:70]
  wire [3:0] drainIdx = _candidateVec_T_1 ? 4'h0 : _drainIdx_T_13; // @[Mux.scala 47:70]
  wire [29:0] inptags_0 = io_in_0_bits_addr[35:6]; // @[Sbuffer.scala 300:7]
  wire [29:0] inptags_1 = io_in_1_bits_addr[35:6]; // @[Sbuffer.scala 300:7]
  wire [32:0] invtags_0 = io_in_0_bits_vaddr[38:6]; // @[Sbuffer.scala 303:7]
  wire [32:0] invtags_1 = io_in_1_bits_vaddr[38:6]; // @[Sbuffer.scala 303:7]
  wire  sameTag = inptags_0 == inptags_1; // @[Sbuffer.scala 375:28]
  wire [32:0] firstWord = io_in_0_bits_addr[35:3]; // @[Sbuffer.scala 306:7]
  wire [32:0] secondWord = io_in_1_bits_addr[35:3]; // @[Sbuffer.scala 306:7]
  wire  sameWord = firstWord == secondWord; // @[Sbuffer.scala 378:28]
  wire  _T_28 = inptags_0 == ptag_14; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_14 = inptags_0 == ptag_14 & _candidateVec_T_57; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T = mergeMask_0_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire  _T_26 = inptags_0 == ptag_13; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_13 = inptags_0 == ptag_13 & _candidateVec_T_53; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_1 = mergeMask_0_13 ? 4'hd : _mergeIdx_T; // @[Mux.scala 47:70]
  wire  _T_24 = inptags_0 == ptag_12; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_12 = inptags_0 == ptag_12 & _candidateVec_T_49; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_2 = mergeMask_0_12 ? 4'hc : _mergeIdx_T_1; // @[Mux.scala 47:70]
  wire  _T_22 = inptags_0 == ptag_11; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_11 = inptags_0 == ptag_11 & _candidateVec_T_45; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_3 = mergeMask_0_11 ? 4'hb : _mergeIdx_T_2; // @[Mux.scala 47:70]
  wire  _T_20 = inptags_0 == ptag_10; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_10 = inptags_0 == ptag_10 & _candidateVec_T_41; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_4 = mergeMask_0_10 ? 4'ha : _mergeIdx_T_3; // @[Mux.scala 47:70]
  wire  _T_18 = inptags_0 == ptag_9; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_9 = inptags_0 == ptag_9 & _candidateVec_T_37; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_5 = mergeMask_0_9 ? 4'h9 : _mergeIdx_T_4; // @[Mux.scala 47:70]
  wire  _T_16 = inptags_0 == ptag_8; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_8 = inptags_0 == ptag_8 & _candidateVec_T_33; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_6 = mergeMask_0_8 ? 4'h8 : _mergeIdx_T_5; // @[Mux.scala 47:70]
  wire  _T_14 = inptags_0 == ptag_7; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_7 = inptags_0 == ptag_7 & _candidateVec_T_29; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_7 = mergeMask_0_7 ? 4'h7 : _mergeIdx_T_6; // @[Mux.scala 47:70]
  wire  _T_12 = inptags_0 == ptag_6; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_6 = inptags_0 == ptag_6 & _candidateVec_T_25; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_8 = mergeMask_0_6 ? 4'h6 : _mergeIdx_T_7; // @[Mux.scala 47:70]
  wire  _T_10 = inptags_0 == ptag_5; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_5 = inptags_0 == ptag_5 & _candidateVec_T_21; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_9 = mergeMask_0_5 ? 4'h5 : _mergeIdx_T_8; // @[Mux.scala 47:70]
  wire  _T_8 = inptags_0 == ptag_4; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_4 = inptags_0 == ptag_4 & _candidateVec_T_17; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_10 = mergeMask_0_4 ? 4'h4 : _mergeIdx_T_9; // @[Mux.scala 47:70]
  wire  _T_6 = inptags_0 == ptag_3; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_3 = inptags_0 == ptag_3 & _candidateVec_T_13; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_11 = mergeMask_0_3 ? 4'h3 : _mergeIdx_T_10; // @[Mux.scala 47:70]
  wire  _T_4 = inptags_0 == ptag_2; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_2 = inptags_0 == ptag_2 & _candidateVec_T_9; // @[Sbuffer.scala 388:30]
  wire  _T_2 = inptags_0 == ptag_1; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_1 = inptags_0 == ptag_1 & _candidateVec_T_5; // @[Sbuffer.scala 388:30]
  wire  _T = inptags_0 == ptag_0; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_0 = inptags_0 == ptag_0 & _candidateVec_T_1; // @[Sbuffer.scala 388:30]
  wire  _T_114 = inptags_1 == ptag_14; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_14 = inptags_1 == ptag_14 & _candidateVec_T_57; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_14 = mergeMask_1_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire  _T_112 = inptags_1 == ptag_13; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_13 = inptags_1 == ptag_13 & _candidateVec_T_53; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_15 = mergeMask_1_13 ? 4'hd : _mergeIdx_T_14; // @[Mux.scala 47:70]
  wire  _T_110 = inptags_1 == ptag_12; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_12 = inptags_1 == ptag_12 & _candidateVec_T_49; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_16 = mergeMask_1_12 ? 4'hc : _mergeIdx_T_15; // @[Mux.scala 47:70]
  wire  _T_108 = inptags_1 == ptag_11; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_11 = inptags_1 == ptag_11 & _candidateVec_T_45; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_17 = mergeMask_1_11 ? 4'hb : _mergeIdx_T_16; // @[Mux.scala 47:70]
  wire  _T_106 = inptags_1 == ptag_10; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_10 = inptags_1 == ptag_10 & _candidateVec_T_41; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_18 = mergeMask_1_10 ? 4'ha : _mergeIdx_T_17; // @[Mux.scala 47:70]
  wire  _T_104 = inptags_1 == ptag_9; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_9 = inptags_1 == ptag_9 & _candidateVec_T_37; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_19 = mergeMask_1_9 ? 4'h9 : _mergeIdx_T_18; // @[Mux.scala 47:70]
  wire  _T_102 = inptags_1 == ptag_8; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_8 = inptags_1 == ptag_8 & _candidateVec_T_33; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_20 = mergeMask_1_8 ? 4'h8 : _mergeIdx_T_19; // @[Mux.scala 47:70]
  wire  _T_100 = inptags_1 == ptag_7; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_7 = inptags_1 == ptag_7 & _candidateVec_T_29; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_21 = mergeMask_1_7 ? 4'h7 : _mergeIdx_T_20; // @[Mux.scala 47:70]
  wire  _T_98 = inptags_1 == ptag_6; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_6 = inptags_1 == ptag_6 & _candidateVec_T_25; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_22 = mergeMask_1_6 ? 4'h6 : _mergeIdx_T_21; // @[Mux.scala 47:70]
  wire  _T_96 = inptags_1 == ptag_5; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_5 = inptags_1 == ptag_5 & _candidateVec_T_21; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_23 = mergeMask_1_5 ? 4'h5 : _mergeIdx_T_22; // @[Mux.scala 47:70]
  wire  _T_94 = inptags_1 == ptag_4; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_4 = inptags_1 == ptag_4 & _candidateVec_T_17; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_24 = mergeMask_1_4 ? 4'h4 : _mergeIdx_T_23; // @[Mux.scala 47:70]
  wire  _T_92 = inptags_1 == ptag_3; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_3 = inptags_1 == ptag_3 & _candidateVec_T_13; // @[Sbuffer.scala 388:30]
  wire [3:0] _mergeIdx_T_25 = mergeMask_1_3 ? 4'h3 : _mergeIdx_T_24; // @[Mux.scala 47:70]
  wire  _T_90 = inptags_1 == ptag_2; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_2 = inptags_1 == ptag_2 & _candidateVec_T_9; // @[Sbuffer.scala 388:30]
  wire  _T_88 = inptags_1 == ptag_1; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_1 = inptags_1 == ptag_1 & _candidateVec_T_5; // @[Sbuffer.scala 388:30]
  wire  _T_86 = inptags_1 == ptag_0; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_0 = inptags_1 == ptag_0 & _candidateVec_T_1; // @[Sbuffer.scala 388:30]
  wire  _T_30 = inptags_0 == ptag_15; // @[Sbuffer.scala 388:18]
  wire  mergeMask_0_15 = inptags_0 == ptag_15 & _candidateVec_T_61; // @[Sbuffer.scala 388:30]
  wire  canMerge_0 = mergeMask_0_0 | mergeMask_0_1 | (mergeMask_0_2 | mergeMask_0_3) | (mergeMask_0_4 | mergeMask_0_5 |
    (mergeMask_0_6 | mergeMask_0_7)) | (mergeMask_0_8 | mergeMask_0_9 | (mergeMask_0_10 | mergeMask_0_11) | (
    mergeMask_0_12 | mergeMask_0_13 | (mergeMask_0_14 | mergeMask_0_15))); // @[ParallelMux.scala 39:55]
  wire  _T_116 = inptags_1 == ptag_15; // @[Sbuffer.scala 388:18]
  wire  mergeMask_1_15 = inptags_1 == ptag_15 & _candidateVec_T_61; // @[Sbuffer.scala 388:30]
  wire  canMerge_1 = mergeMask_1_0 | mergeMask_1_1 | (mergeMask_1_2 | mergeMask_1_3) | (mergeMask_1_4 | mergeMask_1_5 |
    (mergeMask_1_6 | mergeMask_1_7)) | (mergeMask_1_8 | mergeMask_1_9 | (mergeMask_1_10 | mergeMask_1_11) | (
    mergeMask_1_12 | mergeMask_1_13 | (mergeMask_1_14 | mergeMask_1_15))); // @[ParallelMux.scala 39:55]
  wire [7:0] mergeVec_lo = {mergeMask_0_7,mergeMask_0_6,mergeMask_0_5,mergeMask_0_4,mergeMask_0_3,mergeMask_0_2,
    mergeMask_0_1,mergeMask_0_0}; // @[Sbuffer.scala 384:34]
  wire [15:0] mergeVec_0 = {mergeMask_0_15,mergeMask_0_14,mergeMask_0_13,mergeMask_0_12,mergeMask_0_11,mergeMask_0_10,
    mergeMask_0_9,mergeMask_0_8,mergeVec_lo}; // @[Sbuffer.scala 384:34]
  wire [7:0] mergeVec_lo_1 = {mergeMask_1_7,mergeMask_1_6,mergeMask_1_5,mergeMask_1_4,mergeMask_1_3,mergeMask_1_2,
    mergeMask_1_1,mergeMask_1_0}; // @[Sbuffer.scala 384:34]
  wire [15:0] mergeVec_1 = {mergeMask_1_15,mergeMask_1_14,mergeMask_1_13,mergeMask_1_12,mergeMask_1_11,mergeMask_1_10,
    mergeMask_1_9,mergeMask_1_8,mergeVec_lo_1}; // @[Sbuffer.scala 384:34]
  wire  invalidMask_0 = ~stateVec_0_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_1 = ~stateVec_1_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_2 = ~stateVec_2_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_3 = ~stateVec_3_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_4 = ~stateVec_4_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_5 = ~stateVec_5_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_6 = ~stateVec_6_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_7 = ~stateVec_7_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_8 = ~stateVec_8_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_9 = ~stateVec_9_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_10 = ~stateVec_10_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_11 = ~stateVec_11_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_12 = ~stateVec_12_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_13 = ~stateVec_13_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_14 = ~stateVec_14_state_valid; // @[Sbuffer.scala 62:27]
  wire  invalidMask_15 = ~stateVec_15_state_valid; // @[Sbuffer.scala 62:27]
  wire [7:0] evenInvalidMask_lo = {invalidMask_7,invalidMask_6,invalidMask_5,invalidMask_4,invalidMask_3,invalidMask_2,
    invalidMask_1,invalidMask_0}; // @[Sbuffer.scala 398:49]
  wire [15:0] _evenInvalidMask_T = {invalidMask_15,invalidMask_14,invalidMask_13,invalidMask_12,invalidMask_11,
    invalidMask_10,invalidMask_9,invalidMask_8,evenInvalidMask_lo}; // @[Sbuffer.scala 398:49]
  wire [7:0] evenInvalidMask = {_evenInvalidMask_T[14],_evenInvalidMask_T[12],_evenInvalidMask_T[10],_evenInvalidMask_T[
    8],_evenInvalidMask_T[6],_evenInvalidMask_T[4],_evenInvalidMask_T[2],_evenInvalidMask_T[0]}; // @[BitUtils.scala 185:64]
  wire [7:0] oddInvalidMask = {_evenInvalidMask_T[15],_evenInvalidMask_T[13],_evenInvalidMask_T[11],_evenInvalidMask_T[9
    ],_evenInvalidMask_T[7],_evenInvalidMask_T[5],_evenInvalidMask_T[3],_evenInvalidMask_T[1]}; // @[BitUtils.scala 197:66]
  wire  evenRawInsertVec_output_0 = evenInvalidMask[0]; // @[Sbuffer.scala 403:41]
  wire  evenRawInsertVec_output_1 = ~(|evenRawInsertVec_output_0) & evenInvalidMask[1]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_2 = ~(|evenInvalidMask[1:0]) & evenInvalidMask[2]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_3 = ~(|evenInvalidMask[2:0]) & evenInvalidMask[3]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_4 = ~(|evenInvalidMask[3:0]) & evenInvalidMask[4]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_5 = ~(|evenInvalidMask[4:0]) & evenInvalidMask[5]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_6 = ~(|evenInvalidMask[5:0]) & evenInvalidMask[6]; // @[Sbuffer.scala 405:41]
  wire  evenRawInsertVec_output_7 = ~(|evenInvalidMask[6:0]) & evenInvalidMask[7]; // @[Sbuffer.scala 405:41]
  wire [7:0] evenRawInsertVec = {evenRawInsertVec_output_7,evenRawInsertVec_output_6,evenRawInsertVec_output_5,
    evenRawInsertVec_output_4,evenRawInsertVec_output_3,evenRawInsertVec_output_2,evenRawInsertVec_output_1,
    evenRawInsertVec_output_0}; // @[Sbuffer.scala 407:12]
  wire  oddRawInsertVec_output_0 = oddInvalidMask[0]; // @[Sbuffer.scala 403:41]
  wire  oddRawInsertVec_output_1 = ~(|oddRawInsertVec_output_0) & oddInvalidMask[1]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_2 = ~(|oddInvalidMask[1:0]) & oddInvalidMask[2]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_3 = ~(|oddInvalidMask[2:0]) & oddInvalidMask[3]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_4 = ~(|oddInvalidMask[3:0]) & oddInvalidMask[4]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_5 = ~(|oddInvalidMask[4:0]) & oddInvalidMask[5]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_6 = ~(|oddInvalidMask[5:0]) & oddInvalidMask[6]; // @[Sbuffer.scala 405:41]
  wire  oddRawInsertVec_output_7 = ~(|oddInvalidMask[6:0]) & oddInvalidMask[7]; // @[Sbuffer.scala 405:41]
  wire [7:0] oddRawInsertVec = {oddRawInsertVec_output_7,oddRawInsertVec_output_6,oddRawInsertVec_output_5,
    oddRawInsertVec_output_4,oddRawInsertVec_output_3,oddRawInsertVec_output_2,oddRawInsertVec_output_1,
    oddRawInsertVec_output_0}; // @[Sbuffer.scala 407:12]
  wire  f_tail_28 = evenInvalidMask[6] | evenInvalidMask[7]; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_29 = evenInvalidMask[5] | f_tail_28; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_30 = evenInvalidMask[4] | f_tail_29; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_31 = evenInvalidMask[3] | f_tail_30; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_32 = evenInvalidMask[2] | f_tail_31; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_33 = evenInvalidMask[1] | f_tail_32; // @[PriorityMuxDefault.scala 46:46]
  wire  evenCanInsert = evenRawInsertVec_output_0 | f_tail_33; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_34 = oddInvalidMask[6] | oddInvalidMask[7]; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_35 = oddInvalidMask[5] | f_tail_34; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_36 = oddInvalidMask[4] | f_tail_35; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_37 = oddInvalidMask[3] | f_tail_36; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_38 = oddInvalidMask[2] | f_tail_37; // @[PriorityMuxDefault.scala 46:46]
  wire  f_tail_39 = oddInvalidMask[1] | f_tail_38; // @[PriorityMuxDefault.scala 46:46]
  wire  oddCanInsert = oddRawInsertVec_output_0 | f_tail_39; // @[PriorityMuxDefault.scala 46:46]
  wire [7:0] evenInsertVec_lo = {1'h0,evenRawInsertVec[3],1'h0,evenRawInsertVec[2],1'h0,evenRawInsertVec[1],1'h0,
    evenRawInsertVec[0]}; // @[BitUtils.scala 190:9]
  wire [15:0] evenInsertVec = {1'h0,evenRawInsertVec[7],1'h0,evenRawInsertVec[6],1'h0,evenRawInsertVec[5],1'h0,
    evenRawInsertVec[4],evenInsertVec_lo}; // @[BitUtils.scala 190:9]
  wire [7:0] oddInsertVec_lo = {oddRawInsertVec[3],1'h0,oddRawInsertVec[2],1'h0,oddRawInsertVec[1],1'h0,oddRawInsertVec[
    0],1'h0}; // @[BitUtils.scala 202:9]
  wire [15:0] oddInsertVec = {oddRawInsertVec[7],1'h0,oddRawInsertVec[6],1'h0,oddRawInsertVec[5],1'h0,oddRawInsertVec[4]
    ,1'h0,oddInsertVec_lo}; // @[BitUtils.scala 202:9]
  reg  enbufferSelReg; // @[Sbuffer.scala 419:31]
  wire  _enbufferSelReg_T = ~enbufferSelReg; // @[Sbuffer.scala 421:23]
  wire [15:0] firstInsertVec = enbufferSelReg ? evenInsertVec : oddInsertVec; // @[Sbuffer.scala 429:27]
  wire [15:0] _secondInsertVec_T_1 = _enbufferSelReg_T ? evenInsertVec : oddInsertVec; // @[Sbuffer.scala 432:8]
  wire [15:0] secondInsertVec = sameTag ? firstInsertVec : _secondInsertVec_T_1; // @[Sbuffer.scala 430:28]
  wire  _firstCanInsert_T = sbuffer_state != 2'h3; // @[Sbuffer.scala 434:38]
  wire  _firstCanInsert_T_1 = enbufferSelReg ? evenCanInsert : oddCanInsert; // @[Sbuffer.scala 434:64]
  wire  firstCanInsert = sbuffer_state != 2'h3 & _firstCanInsert_T_1; // @[Sbuffer.scala 434:58]
  wire  _secondCanInsert_T_2 = _enbufferSelReg_T ? evenCanInsert : oddCanInsert; // @[Sbuffer.scala 437:8]
  wire  _secondCanInsert_T_3 = sameTag ? firstCanInsert : _secondCanInsert_T_2; // @[Sbuffer.scala 435:65]
  wire  secondCanInsert = _firstCanInsert_T & _secondCanInsert_T_3; // @[Sbuffer.scala 435:59]
  reg  do_uarch_drain_REG; // @[Sbuffer.scala 441:31]
  reg  do_uarch_drain_REG_1; // @[Sbuffer.scala 441:76]
  reg  do_uarch_drain_REG_2; // @[Sbuffer.scala 441:68]
  wire  do_uarch_drain = do_uarch_drain_REG | do_uarch_drain_REG_2; // @[Sbuffer.scala 441:58]
  wire  _dataModule_io_writeReq_0_valid_T = io_in_0_ready & io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [7:0] insertIdx_hi = firstInsertVec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] insertIdx_lo = firstInsertVec[7:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T = |insertIdx_hi; // @[OneHot.scala 32:14]
  wire [7:0] _insertIdx_T_1 = insertIdx_hi | insertIdx_lo; // @[OneHot.scala 32:28]
  wire [3:0] insertIdx_hi_1 = _insertIdx_T_1[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] insertIdx_lo_1 = _insertIdx_T_1[3:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T_2 = |insertIdx_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _insertIdx_T_3 = insertIdx_hi_1 | insertIdx_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] insertIdx_hi_2 = _insertIdx_T_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] insertIdx_lo_2 = _insertIdx_T_3[1:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T_4 = |insertIdx_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _insertIdx_T_5 = insertIdx_hi_2 | insertIdx_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] insertIdx = {_insertIdx_T,_insertIdx_T_2,_insertIdx_T_4,_insertIdx_T_5[1]}; // @[Cat.scala 33:92]
  reg  accessIdx_0_valid_REG; // @[Sbuffer.scala 509:34]
  reg [3:0] accessIdx_0_bits_REG; // @[Sbuffer.scala 510:33]
  wire  _T_248 = invtags_0 != vtag_0; // @[Sbuffer.scala 486:22]
  wire [20:0] _GEN_3 = mergeVec_0[0] ? 21'h0 : cohCount_0; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_4 = mergeVec_0[0] & _T_248; // @[Sbuffer.scala 482:32 440:40]
  wire  _GEN_5 = invtags_0 != vtag_1 | _GEN_4; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_6 = mergeVec_0[1] ? 21'h0 : cohCount_1; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_7 = mergeVec_0[1] ? _GEN_5 : _GEN_4; // @[Sbuffer.scala 482:32]
  wire  _GEN_8 = invtags_0 != vtag_2 | _GEN_7; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_9 = mergeVec_0[2] ? 21'h0 : cohCount_2; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_10 = mergeVec_0[2] ? _GEN_8 : _GEN_7; // @[Sbuffer.scala 482:32]
  wire  _GEN_11 = invtags_0 != vtag_3 | _GEN_10; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_12 = mergeVec_0[3] ? 21'h0 : cohCount_3; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_13 = mergeVec_0[3] ? _GEN_11 : _GEN_10; // @[Sbuffer.scala 482:32]
  wire  _GEN_14 = invtags_0 != vtag_4 | _GEN_13; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_15 = mergeVec_0[4] ? 21'h0 : cohCount_4; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_16 = mergeVec_0[4] ? _GEN_14 : _GEN_13; // @[Sbuffer.scala 482:32]
  wire  _GEN_17 = invtags_0 != vtag_5 | _GEN_16; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_18 = mergeVec_0[5] ? 21'h0 : cohCount_5; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_19 = mergeVec_0[5] ? _GEN_17 : _GEN_16; // @[Sbuffer.scala 482:32]
  wire  _GEN_20 = invtags_0 != vtag_6 | _GEN_19; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_21 = mergeVec_0[6] ? 21'h0 : cohCount_6; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_22 = mergeVec_0[6] ? _GEN_20 : _GEN_19; // @[Sbuffer.scala 482:32]
  wire  _GEN_23 = invtags_0 != vtag_7 | _GEN_22; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_24 = mergeVec_0[7] ? 21'h0 : cohCount_7; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_25 = mergeVec_0[7] ? _GEN_23 : _GEN_22; // @[Sbuffer.scala 482:32]
  wire  _GEN_26 = invtags_0 != vtag_8 | _GEN_25; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_27 = mergeVec_0[8] ? 21'h0 : cohCount_8; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_28 = mergeVec_0[8] ? _GEN_26 : _GEN_25; // @[Sbuffer.scala 482:32]
  wire  _GEN_29 = invtags_0 != vtag_9 | _GEN_28; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_30 = mergeVec_0[9] ? 21'h0 : cohCount_9; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_31 = mergeVec_0[9] ? _GEN_29 : _GEN_28; // @[Sbuffer.scala 482:32]
  wire  _GEN_32 = invtags_0 != vtag_10 | _GEN_31; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_33 = mergeVec_0[10] ? 21'h0 : cohCount_10; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_34 = mergeVec_0[10] ? _GEN_32 : _GEN_31; // @[Sbuffer.scala 482:32]
  wire  _GEN_35 = invtags_0 != vtag_11 | _GEN_34; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_36 = mergeVec_0[11] ? 21'h0 : cohCount_11; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_37 = mergeVec_0[11] ? _GEN_35 : _GEN_34; // @[Sbuffer.scala 482:32]
  wire  _GEN_38 = invtags_0 != vtag_12 | _GEN_37; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_39 = mergeVec_0[12] ? 21'h0 : cohCount_12; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_40 = mergeVec_0[12] ? _GEN_38 : _GEN_37; // @[Sbuffer.scala 482:32]
  wire  _GEN_41 = invtags_0 != vtag_13 | _GEN_40; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_42 = mergeVec_0[13] ? 21'h0 : cohCount_13; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_43 = mergeVec_0[13] ? _GEN_41 : _GEN_40; // @[Sbuffer.scala 482:32]
  wire  _GEN_44 = invtags_0 != vtag_14 | _GEN_43; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_45 = mergeVec_0[14] ? 21'h0 : cohCount_14; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_46 = mergeVec_0[14] ? _GEN_44 : _GEN_43; // @[Sbuffer.scala 482:32]
  wire  _GEN_47 = invtags_0 != vtag_15 | _GEN_46; // @[Sbuffer.scala 486:42 493:34]
  wire [20:0] _GEN_48 = mergeVec_0[15] ? 21'h0 : cohCount_15; // @[Sbuffer.scala 281:25 482:32 483:28]
  wire  _GEN_49 = mergeVec_0[15] ? _GEN_47 : _GEN_46; // @[Sbuffer.scala 482:32]
  wire  _sameBlockInflightMask_mask_T_1 = stateVec_0_state_inflight & _T; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_3 = stateVec_1_state_inflight & _T_2; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_5 = stateVec_2_state_inflight & _T_4; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_7 = stateVec_3_state_inflight & _T_6; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_9 = stateVec_4_state_inflight & _T_8; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_11 = stateVec_5_state_inflight & _T_10; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_13 = stateVec_6_state_inflight & _T_12; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_15 = stateVec_7_state_inflight & _T_14; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_17 = stateVec_8_state_inflight & _T_16; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_19 = stateVec_9_state_inflight & _T_18; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_21 = stateVec_10_state_inflight & _T_20; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_23 = stateVec_11_state_inflight & _T_22; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_25 = stateVec_12_state_inflight & _T_24; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_27 = stateVec_13_state_inflight & _T_26; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_29 = stateVec_14_state_inflight & _T_28; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_31 = stateVec_15_state_inflight & _T_30; // @[Sbuffer.scala 599:54]
  wire [7:0] sameBlockInflightMask_mask_lo = {_sameBlockInflightMask_mask_T_15,_sameBlockInflightMask_mask_T_13,
    _sameBlockInflightMask_mask_T_11,_sameBlockInflightMask_mask_T_9,_sameBlockInflightMask_mask_T_7,
    _sameBlockInflightMask_mask_T_5,_sameBlockInflightMask_mask_T_3,_sameBlockInflightMask_mask_T_1}; // @[Sbuffer.scala 599:79]
  wire [15:0] sameBlockInflightMask = {_sameBlockInflightMask_mask_T_31,_sameBlockInflightMask_mask_T_29,
    _sameBlockInflightMask_mask_T_27,_sameBlockInflightMask_mask_T_25,_sameBlockInflightMask_mask_T_23,
    _sameBlockInflightMask_mask_T_21,_sameBlockInflightMask_mask_T_19,_sameBlockInflightMask_mask_T_17,
    sameBlockInflightMask_mask_lo}; // @[Sbuffer.scala 599:79]
  wire  _stateVec_0_w_sameblock_inflight_T = |sameBlockInflightMask; // @[Sbuffer.scala 460:74]
  wire [15:0] _GEN_50 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_0; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_51 = firstInsertVec[0] | stateVec_0_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_52 = firstInsertVec[0] ? |sameBlockInflightMask : stateVec_0_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_53 = firstInsertVec[0] ? _GEN_50 : waitInflightMask_0; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_54 = firstInsertVec[0] ? 21'h0 : cohCount_0; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_55 = firstInsertVec[0] ? inptags_0 : ptag_0; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_56 = firstInsertVec[0] ? invtags_0 : vtag_0; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_57 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_1; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_58 = firstInsertVec[1] | stateVec_1_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_59 = firstInsertVec[1] ? |sameBlockInflightMask : stateVec_1_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_60 = firstInsertVec[1] ? _GEN_57 : waitInflightMask_1; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_61 = firstInsertVec[1] ? 21'h0 : cohCount_1; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_62 = firstInsertVec[1] ? inptags_0 : ptag_1; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_63 = firstInsertVec[1] ? invtags_0 : vtag_1; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_64 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_2; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_65 = firstInsertVec[2] | stateVec_2_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_66 = firstInsertVec[2] ? |sameBlockInflightMask : stateVec_2_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_67 = firstInsertVec[2] ? _GEN_64 : waitInflightMask_2; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_68 = firstInsertVec[2] ? 21'h0 : cohCount_2; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_69 = firstInsertVec[2] ? inptags_0 : ptag_2; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_70 = firstInsertVec[2] ? invtags_0 : vtag_2; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_71 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_3; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_72 = firstInsertVec[3] | stateVec_3_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_73 = firstInsertVec[3] ? |sameBlockInflightMask : stateVec_3_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_74 = firstInsertVec[3] ? _GEN_71 : waitInflightMask_3; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_75 = firstInsertVec[3] ? 21'h0 : cohCount_3; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_76 = firstInsertVec[3] ? inptags_0 : ptag_3; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_77 = firstInsertVec[3] ? invtags_0 : vtag_3; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_78 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_4; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_79 = firstInsertVec[4] | stateVec_4_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_80 = firstInsertVec[4] ? |sameBlockInflightMask : stateVec_4_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_81 = firstInsertVec[4] ? _GEN_78 : waitInflightMask_4; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_82 = firstInsertVec[4] ? 21'h0 : cohCount_4; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_83 = firstInsertVec[4] ? inptags_0 : ptag_4; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_84 = firstInsertVec[4] ? invtags_0 : vtag_4; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_85 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_5; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_86 = firstInsertVec[5] | stateVec_5_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_87 = firstInsertVec[5] ? |sameBlockInflightMask : stateVec_5_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_88 = firstInsertVec[5] ? _GEN_85 : waitInflightMask_5; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_89 = firstInsertVec[5] ? 21'h0 : cohCount_5; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_90 = firstInsertVec[5] ? inptags_0 : ptag_5; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_91 = firstInsertVec[5] ? invtags_0 : vtag_5; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_92 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_6; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_93 = firstInsertVec[6] | stateVec_6_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_94 = firstInsertVec[6] ? |sameBlockInflightMask : stateVec_6_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_95 = firstInsertVec[6] ? _GEN_92 : waitInflightMask_6; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_96 = firstInsertVec[6] ? 21'h0 : cohCount_6; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_97 = firstInsertVec[6] ? inptags_0 : ptag_6; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_98 = firstInsertVec[6] ? invtags_0 : vtag_6; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_99 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_7; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_100 = firstInsertVec[7] | stateVec_7_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_101 = firstInsertVec[7] ? |sameBlockInflightMask : stateVec_7_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_102 = firstInsertVec[7] ? _GEN_99 : waitInflightMask_7; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_103 = firstInsertVec[7] ? 21'h0 : cohCount_7; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_104 = firstInsertVec[7] ? inptags_0 : ptag_7; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_105 = firstInsertVec[7] ? invtags_0 : vtag_7; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_106 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_8; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_107 = firstInsertVec[8] | stateVec_8_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_108 = firstInsertVec[8] ? |sameBlockInflightMask : stateVec_8_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_109 = firstInsertVec[8] ? _GEN_106 : waitInflightMask_8; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_110 = firstInsertVec[8] ? 21'h0 : cohCount_8; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_111 = firstInsertVec[8] ? inptags_0 : ptag_8; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_112 = firstInsertVec[8] ? invtags_0 : vtag_8; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_113 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_9; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_114 = firstInsertVec[9] | stateVec_9_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_115 = firstInsertVec[9] ? |sameBlockInflightMask : stateVec_9_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_116 = firstInsertVec[9] ? _GEN_113 : waitInflightMask_9; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_117 = firstInsertVec[9] ? 21'h0 : cohCount_9; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_118 = firstInsertVec[9] ? inptags_0 : ptag_9; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_119 = firstInsertVec[9] ? invtags_0 : vtag_9; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_120 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_10; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_121 = firstInsertVec[10] | stateVec_10_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_122 = firstInsertVec[10] ? |sameBlockInflightMask : stateVec_10_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_123 = firstInsertVec[10] ? _GEN_120 : waitInflightMask_10; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_124 = firstInsertVec[10] ? 21'h0 : cohCount_10; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_125 = firstInsertVec[10] ? inptags_0 : ptag_10; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_126 = firstInsertVec[10] ? invtags_0 : vtag_10; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_127 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_11; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_128 = firstInsertVec[11] | stateVec_11_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_129 = firstInsertVec[11] ? |sameBlockInflightMask : stateVec_11_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_130 = firstInsertVec[11] ? _GEN_127 : waitInflightMask_11; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_131 = firstInsertVec[11] ? 21'h0 : cohCount_11; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_132 = firstInsertVec[11] ? inptags_0 : ptag_11; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_133 = firstInsertVec[11] ? invtags_0 : vtag_11; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_134 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_12; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_135 = firstInsertVec[12] | stateVec_12_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_136 = firstInsertVec[12] ? |sameBlockInflightMask : stateVec_12_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_137 = firstInsertVec[12] ? _GEN_134 : waitInflightMask_12; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_138 = firstInsertVec[12] ? 21'h0 : cohCount_12; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_139 = firstInsertVec[12] ? inptags_0 : ptag_12; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_140 = firstInsertVec[12] ? invtags_0 : vtag_12; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_141 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_13; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_142 = firstInsertVec[13] | stateVec_13_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_143 = firstInsertVec[13] ? |sameBlockInflightMask : stateVec_13_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_144 = firstInsertVec[13] ? _GEN_141 : waitInflightMask_13; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_145 = firstInsertVec[13] ? 21'h0 : cohCount_13; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_146 = firstInsertVec[13] ? inptags_0 : ptag_13; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_147 = firstInsertVec[13] ? invtags_0 : vtag_13; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_148 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_14; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_149 = firstInsertVec[14] | stateVec_14_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_150 = firstInsertVec[14] ? |sameBlockInflightMask : stateVec_14_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_151 = firstInsertVec[14] ? _GEN_148 : waitInflightMask_14; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_152 = firstInsertVec[14] ? 21'h0 : cohCount_14; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_153 = firstInsertVec[14] ? inptags_0 : ptag_14; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_154 = firstInsertVec[14] ? invtags_0 : vtag_14; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [15:0] _GEN_155 = _stateVec_0_w_sameblock_inflight_T ? sameBlockInflightMask : waitInflightMask_15; // @[Sbuffer.scala 277:29 461:40 462:38]
  wire  _GEN_156 = firstInsertVec[15] | stateVec_15_state_valid; // @[Sbuffer.scala 280:25 458:32 459:40]
  wire  _GEN_157 = firstInsertVec[15] ? |sameBlockInflightMask : stateVec_15_w_sameblock_inflight; // @[Sbuffer.scala 280:25 458:32 460:49]
  wire [15:0] _GEN_158 = firstInsertVec[15] ? _GEN_155 : waitInflightMask_15; // @[Sbuffer.scala 277:29 458:32]
  wire [20:0] _GEN_159 = firstInsertVec[15] ? 21'h0 : cohCount_15; // @[Sbuffer.scala 281:25 458:32 464:28]
  wire [29:0] _GEN_160 = firstInsertVec[15] ? inptags_0 : ptag_15; // @[Sbuffer.scala 274:17 458:32 466:24]
  wire [32:0] _GEN_161 = firstInsertVec[15] ? invtags_0 : vtag_15; // @[Sbuffer.scala 275:17 458:32 467:24]
  wire [20:0] _GEN_163 = canMerge_0 ? _GEN_3 : _GEN_54; // @[Sbuffer.scala 512:24]
  wire  _GEN_164 = canMerge_0 & _GEN_49; // @[Sbuffer.scala 512:24 440:40]
  wire [20:0] _GEN_165 = canMerge_0 ? _GEN_6 : _GEN_61; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_166 = canMerge_0 ? _GEN_9 : _GEN_68; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_167 = canMerge_0 ? _GEN_12 : _GEN_75; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_168 = canMerge_0 ? _GEN_15 : _GEN_82; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_169 = canMerge_0 ? _GEN_18 : _GEN_89; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_170 = canMerge_0 ? _GEN_21 : _GEN_96; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_171 = canMerge_0 ? _GEN_24 : _GEN_103; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_172 = canMerge_0 ? _GEN_27 : _GEN_110; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_173 = canMerge_0 ? _GEN_30 : _GEN_117; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_174 = canMerge_0 ? _GEN_33 : _GEN_124; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_175 = canMerge_0 ? _GEN_36 : _GEN_131; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_176 = canMerge_0 ? _GEN_39 : _GEN_138; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_177 = canMerge_0 ? _GEN_42 : _GEN_145; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_178 = canMerge_0 ? _GEN_45 : _GEN_152; // @[Sbuffer.scala 512:24]
  wire [20:0] _GEN_179 = canMerge_0 ? _GEN_48 : _GEN_159; // @[Sbuffer.scala 512:24]
  wire  _GEN_180 = canMerge_0 ? stateVec_0_state_valid : _GEN_51; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_181 = canMerge_0 ? stateVec_0_w_sameblock_inflight : _GEN_52; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_182 = canMerge_0 ? waitInflightMask_0 : _GEN_53; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_183 = canMerge_0 ? ptag_0 : _GEN_55; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_184 = canMerge_0 ? vtag_0 : _GEN_56; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_185 = canMerge_0 ? stateVec_1_state_valid : _GEN_58; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_186 = canMerge_0 ? stateVec_1_w_sameblock_inflight : _GEN_59; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_187 = canMerge_0 ? waitInflightMask_1 : _GEN_60; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_188 = canMerge_0 ? ptag_1 : _GEN_62; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_189 = canMerge_0 ? vtag_1 : _GEN_63; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_190 = canMerge_0 ? stateVec_2_state_valid : _GEN_65; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_191 = canMerge_0 ? stateVec_2_w_sameblock_inflight : _GEN_66; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_192 = canMerge_0 ? waitInflightMask_2 : _GEN_67; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_193 = canMerge_0 ? ptag_2 : _GEN_69; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_194 = canMerge_0 ? vtag_2 : _GEN_70; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_195 = canMerge_0 ? stateVec_3_state_valid : _GEN_72; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_196 = canMerge_0 ? stateVec_3_w_sameblock_inflight : _GEN_73; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_197 = canMerge_0 ? waitInflightMask_3 : _GEN_74; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_198 = canMerge_0 ? ptag_3 : _GEN_76; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_199 = canMerge_0 ? vtag_3 : _GEN_77; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_200 = canMerge_0 ? stateVec_4_state_valid : _GEN_79; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_201 = canMerge_0 ? stateVec_4_w_sameblock_inflight : _GEN_80; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_202 = canMerge_0 ? waitInflightMask_4 : _GEN_81; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_203 = canMerge_0 ? ptag_4 : _GEN_83; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_204 = canMerge_0 ? vtag_4 : _GEN_84; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_205 = canMerge_0 ? stateVec_5_state_valid : _GEN_86; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_206 = canMerge_0 ? stateVec_5_w_sameblock_inflight : _GEN_87; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_207 = canMerge_0 ? waitInflightMask_5 : _GEN_88; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_208 = canMerge_0 ? ptag_5 : _GEN_90; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_209 = canMerge_0 ? vtag_5 : _GEN_91; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_210 = canMerge_0 ? stateVec_6_state_valid : _GEN_93; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_211 = canMerge_0 ? stateVec_6_w_sameblock_inflight : _GEN_94; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_212 = canMerge_0 ? waitInflightMask_6 : _GEN_95; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_213 = canMerge_0 ? ptag_6 : _GEN_97; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_214 = canMerge_0 ? vtag_6 : _GEN_98; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_215 = canMerge_0 ? stateVec_7_state_valid : _GEN_100; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_216 = canMerge_0 ? stateVec_7_w_sameblock_inflight : _GEN_101; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_217 = canMerge_0 ? waitInflightMask_7 : _GEN_102; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_218 = canMerge_0 ? ptag_7 : _GEN_104; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_219 = canMerge_0 ? vtag_7 : _GEN_105; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_220 = canMerge_0 ? stateVec_8_state_valid : _GEN_107; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_221 = canMerge_0 ? stateVec_8_w_sameblock_inflight : _GEN_108; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_222 = canMerge_0 ? waitInflightMask_8 : _GEN_109; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_223 = canMerge_0 ? ptag_8 : _GEN_111; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_224 = canMerge_0 ? vtag_8 : _GEN_112; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_225 = canMerge_0 ? stateVec_9_state_valid : _GEN_114; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_226 = canMerge_0 ? stateVec_9_w_sameblock_inflight : _GEN_115; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_227 = canMerge_0 ? waitInflightMask_9 : _GEN_116; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_228 = canMerge_0 ? ptag_9 : _GEN_118; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_229 = canMerge_0 ? vtag_9 : _GEN_119; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_230 = canMerge_0 ? stateVec_10_state_valid : _GEN_121; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_231 = canMerge_0 ? stateVec_10_w_sameblock_inflight : _GEN_122; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_232 = canMerge_0 ? waitInflightMask_10 : _GEN_123; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_233 = canMerge_0 ? ptag_10 : _GEN_125; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_234 = canMerge_0 ? vtag_10 : _GEN_126; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_235 = canMerge_0 ? stateVec_11_state_valid : _GEN_128; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_236 = canMerge_0 ? stateVec_11_w_sameblock_inflight : _GEN_129; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_237 = canMerge_0 ? waitInflightMask_11 : _GEN_130; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_238 = canMerge_0 ? ptag_11 : _GEN_132; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_239 = canMerge_0 ? vtag_11 : _GEN_133; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_240 = canMerge_0 ? stateVec_12_state_valid : _GEN_135; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_241 = canMerge_0 ? stateVec_12_w_sameblock_inflight : _GEN_136; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_242 = canMerge_0 ? waitInflightMask_12 : _GEN_137; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_243 = canMerge_0 ? ptag_12 : _GEN_139; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_244 = canMerge_0 ? vtag_12 : _GEN_140; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_245 = canMerge_0 ? stateVec_13_state_valid : _GEN_142; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_246 = canMerge_0 ? stateVec_13_w_sameblock_inflight : _GEN_143; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_247 = canMerge_0 ? waitInflightMask_13 : _GEN_144; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_248 = canMerge_0 ? ptag_13 : _GEN_146; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_249 = canMerge_0 ? vtag_13 : _GEN_147; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_250 = canMerge_0 ? stateVec_14_state_valid : _GEN_149; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_251 = canMerge_0 ? stateVec_14_w_sameblock_inflight : _GEN_150; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_252 = canMerge_0 ? waitInflightMask_14 : _GEN_151; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_253 = canMerge_0 ? ptag_14 : _GEN_153; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_254 = canMerge_0 ? vtag_14 : _GEN_154; // @[Sbuffer.scala 275:17 512:24]
  wire  _GEN_255 = canMerge_0 ? stateVec_15_state_valid : _GEN_156; // @[Sbuffer.scala 512:24 280:25]
  wire  _GEN_256 = canMerge_0 ? stateVec_15_w_sameblock_inflight : _GEN_157; // @[Sbuffer.scala 512:24 280:25]
  wire [15:0] _GEN_257 = canMerge_0 ? waitInflightMask_15 : _GEN_158; // @[Sbuffer.scala 512:24 277:29]
  wire [29:0] _GEN_258 = canMerge_0 ? ptag_15 : _GEN_160; // @[Sbuffer.scala 274:17 512:24]
  wire [32:0] _GEN_259 = canMerge_0 ? vtag_15 : _GEN_161; // @[Sbuffer.scala 275:17 512:24]
  wire [20:0] _GEN_261 = _dataModule_io_writeReq_0_valid_T ? _GEN_163 : cohCount_0; // @[Sbuffer.scala 511:20 281:25]
  wire  _GEN_262 = _dataModule_io_writeReq_0_valid_T & _GEN_164; // @[Sbuffer.scala 511:20 440:40]
  wire [20:0] _GEN_263 = _dataModule_io_writeReq_0_valid_T ? _GEN_165 : cohCount_1; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_264 = _dataModule_io_writeReq_0_valid_T ? _GEN_166 : cohCount_2; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_265 = _dataModule_io_writeReq_0_valid_T ? _GEN_167 : cohCount_3; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_266 = _dataModule_io_writeReq_0_valid_T ? _GEN_168 : cohCount_4; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_267 = _dataModule_io_writeReq_0_valid_T ? _GEN_169 : cohCount_5; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_268 = _dataModule_io_writeReq_0_valid_T ? _GEN_170 : cohCount_6; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_269 = _dataModule_io_writeReq_0_valid_T ? _GEN_171 : cohCount_7; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_270 = _dataModule_io_writeReq_0_valid_T ? _GEN_172 : cohCount_8; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_271 = _dataModule_io_writeReq_0_valid_T ? _GEN_173 : cohCount_9; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_272 = _dataModule_io_writeReq_0_valid_T ? _GEN_174 : cohCount_10; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_273 = _dataModule_io_writeReq_0_valid_T ? _GEN_175 : cohCount_11; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_274 = _dataModule_io_writeReq_0_valid_T ? _GEN_176 : cohCount_12; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_275 = _dataModule_io_writeReq_0_valid_T ? _GEN_177 : cohCount_13; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_276 = _dataModule_io_writeReq_0_valid_T ? _GEN_178 : cohCount_14; // @[Sbuffer.scala 511:20 281:25]
  wire [20:0] _GEN_277 = _dataModule_io_writeReq_0_valid_T ? _GEN_179 : cohCount_15; // @[Sbuffer.scala 511:20 281:25]
  wire  _GEN_278 = _dataModule_io_writeReq_0_valid_T ? _GEN_180 : stateVec_0_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_279 = _dataModule_io_writeReq_0_valid_T ? _GEN_181 : stateVec_0_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_280 = _dataModule_io_writeReq_0_valid_T ? _GEN_182 : waitInflightMask_0; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_281 = _dataModule_io_writeReq_0_valid_T ? _GEN_183 : ptag_0; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_282 = _dataModule_io_writeReq_0_valid_T ? _GEN_184 : vtag_0; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_283 = _dataModule_io_writeReq_0_valid_T ? _GEN_185 : stateVec_1_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_284 = _dataModule_io_writeReq_0_valid_T ? _GEN_186 : stateVec_1_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_285 = _dataModule_io_writeReq_0_valid_T ? _GEN_187 : waitInflightMask_1; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_286 = _dataModule_io_writeReq_0_valid_T ? _GEN_188 : ptag_1; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_287 = _dataModule_io_writeReq_0_valid_T ? _GEN_189 : vtag_1; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_288 = _dataModule_io_writeReq_0_valid_T ? _GEN_190 : stateVec_2_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_289 = _dataModule_io_writeReq_0_valid_T ? _GEN_191 : stateVec_2_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_290 = _dataModule_io_writeReq_0_valid_T ? _GEN_192 : waitInflightMask_2; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_291 = _dataModule_io_writeReq_0_valid_T ? _GEN_193 : ptag_2; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_292 = _dataModule_io_writeReq_0_valid_T ? _GEN_194 : vtag_2; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_293 = _dataModule_io_writeReq_0_valid_T ? _GEN_195 : stateVec_3_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_294 = _dataModule_io_writeReq_0_valid_T ? _GEN_196 : stateVec_3_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_295 = _dataModule_io_writeReq_0_valid_T ? _GEN_197 : waitInflightMask_3; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_296 = _dataModule_io_writeReq_0_valid_T ? _GEN_198 : ptag_3; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_297 = _dataModule_io_writeReq_0_valid_T ? _GEN_199 : vtag_3; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_298 = _dataModule_io_writeReq_0_valid_T ? _GEN_200 : stateVec_4_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_299 = _dataModule_io_writeReq_0_valid_T ? _GEN_201 : stateVec_4_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_300 = _dataModule_io_writeReq_0_valid_T ? _GEN_202 : waitInflightMask_4; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_301 = _dataModule_io_writeReq_0_valid_T ? _GEN_203 : ptag_4; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_302 = _dataModule_io_writeReq_0_valid_T ? _GEN_204 : vtag_4; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_303 = _dataModule_io_writeReq_0_valid_T ? _GEN_205 : stateVec_5_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_304 = _dataModule_io_writeReq_0_valid_T ? _GEN_206 : stateVec_5_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_305 = _dataModule_io_writeReq_0_valid_T ? _GEN_207 : waitInflightMask_5; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_306 = _dataModule_io_writeReq_0_valid_T ? _GEN_208 : ptag_5; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_307 = _dataModule_io_writeReq_0_valid_T ? _GEN_209 : vtag_5; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_308 = _dataModule_io_writeReq_0_valid_T ? _GEN_210 : stateVec_6_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_309 = _dataModule_io_writeReq_0_valid_T ? _GEN_211 : stateVec_6_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_310 = _dataModule_io_writeReq_0_valid_T ? _GEN_212 : waitInflightMask_6; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_311 = _dataModule_io_writeReq_0_valid_T ? _GEN_213 : ptag_6; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_312 = _dataModule_io_writeReq_0_valid_T ? _GEN_214 : vtag_6; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_313 = _dataModule_io_writeReq_0_valid_T ? _GEN_215 : stateVec_7_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_314 = _dataModule_io_writeReq_0_valid_T ? _GEN_216 : stateVec_7_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_315 = _dataModule_io_writeReq_0_valid_T ? _GEN_217 : waitInflightMask_7; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_316 = _dataModule_io_writeReq_0_valid_T ? _GEN_218 : ptag_7; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_317 = _dataModule_io_writeReq_0_valid_T ? _GEN_219 : vtag_7; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_318 = _dataModule_io_writeReq_0_valid_T ? _GEN_220 : stateVec_8_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_319 = _dataModule_io_writeReq_0_valid_T ? _GEN_221 : stateVec_8_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_320 = _dataModule_io_writeReq_0_valid_T ? _GEN_222 : waitInflightMask_8; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_321 = _dataModule_io_writeReq_0_valid_T ? _GEN_223 : ptag_8; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_322 = _dataModule_io_writeReq_0_valid_T ? _GEN_224 : vtag_8; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_323 = _dataModule_io_writeReq_0_valid_T ? _GEN_225 : stateVec_9_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_324 = _dataModule_io_writeReq_0_valid_T ? _GEN_226 : stateVec_9_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_325 = _dataModule_io_writeReq_0_valid_T ? _GEN_227 : waitInflightMask_9; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_326 = _dataModule_io_writeReq_0_valid_T ? _GEN_228 : ptag_9; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_327 = _dataModule_io_writeReq_0_valid_T ? _GEN_229 : vtag_9; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_328 = _dataModule_io_writeReq_0_valid_T ? _GEN_230 : stateVec_10_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_329 = _dataModule_io_writeReq_0_valid_T ? _GEN_231 : stateVec_10_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_330 = _dataModule_io_writeReq_0_valid_T ? _GEN_232 : waitInflightMask_10; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_331 = _dataModule_io_writeReq_0_valid_T ? _GEN_233 : ptag_10; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_332 = _dataModule_io_writeReq_0_valid_T ? _GEN_234 : vtag_10; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_333 = _dataModule_io_writeReq_0_valid_T ? _GEN_235 : stateVec_11_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_334 = _dataModule_io_writeReq_0_valid_T ? _GEN_236 : stateVec_11_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_335 = _dataModule_io_writeReq_0_valid_T ? _GEN_237 : waitInflightMask_11; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_336 = _dataModule_io_writeReq_0_valid_T ? _GEN_238 : ptag_11; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_337 = _dataModule_io_writeReq_0_valid_T ? _GEN_239 : vtag_11; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_338 = _dataModule_io_writeReq_0_valid_T ? _GEN_240 : stateVec_12_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_339 = _dataModule_io_writeReq_0_valid_T ? _GEN_241 : stateVec_12_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_340 = _dataModule_io_writeReq_0_valid_T ? _GEN_242 : waitInflightMask_12; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_341 = _dataModule_io_writeReq_0_valid_T ? _GEN_243 : ptag_12; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_342 = _dataModule_io_writeReq_0_valid_T ? _GEN_244 : vtag_12; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_343 = _dataModule_io_writeReq_0_valid_T ? _GEN_245 : stateVec_13_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_344 = _dataModule_io_writeReq_0_valid_T ? _GEN_246 : stateVec_13_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_345 = _dataModule_io_writeReq_0_valid_T ? _GEN_247 : waitInflightMask_13; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_346 = _dataModule_io_writeReq_0_valid_T ? _GEN_248 : ptag_13; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_347 = _dataModule_io_writeReq_0_valid_T ? _GEN_249 : vtag_13; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_348 = _dataModule_io_writeReq_0_valid_T ? _GEN_250 : stateVec_14_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_349 = _dataModule_io_writeReq_0_valid_T ? _GEN_251 : stateVec_14_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_350 = _dataModule_io_writeReq_0_valid_T ? _GEN_252 : waitInflightMask_14; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_351 = _dataModule_io_writeReq_0_valid_T ? _GEN_253 : ptag_14; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_352 = _dataModule_io_writeReq_0_valid_T ? _GEN_254 : vtag_14; // @[Sbuffer.scala 275:17 511:20]
  wire  _GEN_353 = _dataModule_io_writeReq_0_valid_T ? _GEN_255 : stateVec_15_state_valid; // @[Sbuffer.scala 511:20 280:25]
  wire  _GEN_354 = _dataModule_io_writeReq_0_valid_T ? _GEN_256 : stateVec_15_w_sameblock_inflight; // @[Sbuffer.scala 511:20 280:25]
  wire [15:0] _GEN_355 = _dataModule_io_writeReq_0_valid_T ? _GEN_257 : waitInflightMask_15; // @[Sbuffer.scala 511:20 277:29]
  wire [29:0] _GEN_356 = _dataModule_io_writeReq_0_valid_T ? _GEN_258 : ptag_15; // @[Sbuffer.scala 274:17 511:20]
  wire [32:0] _GEN_357 = _dataModule_io_writeReq_0_valid_T ? _GEN_259 : vtag_15; // @[Sbuffer.scala 275:17 511:20]
  wire  _dataModule_io_writeReq_1_valid_T = io_in_1_ready & io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [7:0] insertIdx_hi_3 = secondInsertVec[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] insertIdx_lo_3 = secondInsertVec[7:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T_9 = |insertIdx_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _insertIdx_T_10 = insertIdx_hi_3 | insertIdx_lo_3; // @[OneHot.scala 32:28]
  wire [3:0] insertIdx_hi_4 = _insertIdx_T_10[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] insertIdx_lo_4 = _insertIdx_T_10[3:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T_11 = |insertIdx_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _insertIdx_T_12 = insertIdx_hi_4 | insertIdx_lo_4; // @[OneHot.scala 32:28]
  wire [1:0] insertIdx_hi_5 = _insertIdx_T_12[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] insertIdx_lo_5 = _insertIdx_T_12[1:0]; // @[OneHot.scala 31:18]
  wire  _insertIdx_T_13 = |insertIdx_hi_5; // @[OneHot.scala 32:14]
  wire [1:0] _insertIdx_T_14 = insertIdx_hi_5 | insertIdx_lo_5; // @[OneHot.scala 32:28]
  wire [3:0] insertIdx_1 = {_insertIdx_T_9,_insertIdx_T_11,_insertIdx_T_13,_insertIdx_T_14[1]}; // @[Cat.scala 33:92]
  reg  accessIdx_1_valid_REG; // @[Sbuffer.scala 509:34]
  reg [3:0] accessIdx_1_bits_REG; // @[Sbuffer.scala 510:33]
  wire  _GEN_358 = invtags_1 != vtag_0 | _GEN_262; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_360 = mergeVec_1[0] ? _GEN_358 : _GEN_262; // @[Sbuffer.scala 482:32]
  wire  _GEN_361 = invtags_1 != vtag_1 | _GEN_360; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_363 = mergeVec_1[1] ? _GEN_361 : _GEN_360; // @[Sbuffer.scala 482:32]
  wire  _GEN_364 = invtags_1 != vtag_2 | _GEN_363; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_366 = mergeVec_1[2] ? _GEN_364 : _GEN_363; // @[Sbuffer.scala 482:32]
  wire  _GEN_367 = invtags_1 != vtag_3 | _GEN_366; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_369 = mergeVec_1[3] ? _GEN_367 : _GEN_366; // @[Sbuffer.scala 482:32]
  wire  _GEN_370 = invtags_1 != vtag_4 | _GEN_369; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_372 = mergeVec_1[4] ? _GEN_370 : _GEN_369; // @[Sbuffer.scala 482:32]
  wire  _GEN_373 = invtags_1 != vtag_5 | _GEN_372; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_375 = mergeVec_1[5] ? _GEN_373 : _GEN_372; // @[Sbuffer.scala 482:32]
  wire  _GEN_376 = invtags_1 != vtag_6 | _GEN_375; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_378 = mergeVec_1[6] ? _GEN_376 : _GEN_375; // @[Sbuffer.scala 482:32]
  wire  _GEN_379 = invtags_1 != vtag_7 | _GEN_378; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_381 = mergeVec_1[7] ? _GEN_379 : _GEN_378; // @[Sbuffer.scala 482:32]
  wire  _GEN_382 = invtags_1 != vtag_8 | _GEN_381; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_384 = mergeVec_1[8] ? _GEN_382 : _GEN_381; // @[Sbuffer.scala 482:32]
  wire  _GEN_385 = invtags_1 != vtag_9 | _GEN_384; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_387 = mergeVec_1[9] ? _GEN_385 : _GEN_384; // @[Sbuffer.scala 482:32]
  wire  _GEN_388 = invtags_1 != vtag_10 | _GEN_387; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_390 = mergeVec_1[10] ? _GEN_388 : _GEN_387; // @[Sbuffer.scala 482:32]
  wire  _GEN_391 = invtags_1 != vtag_11 | _GEN_390; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_393 = mergeVec_1[11] ? _GEN_391 : _GEN_390; // @[Sbuffer.scala 482:32]
  wire  _GEN_394 = invtags_1 != vtag_12 | _GEN_393; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_396 = mergeVec_1[12] ? _GEN_394 : _GEN_393; // @[Sbuffer.scala 482:32]
  wire  _GEN_397 = invtags_1 != vtag_13 | _GEN_396; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_399 = mergeVec_1[13] ? _GEN_397 : _GEN_396; // @[Sbuffer.scala 482:32]
  wire  _GEN_400 = invtags_1 != vtag_14 | _GEN_399; // @[Sbuffer.scala 486:42 493:34]
  wire  _GEN_402 = mergeVec_1[14] ? _GEN_400 : _GEN_399; // @[Sbuffer.scala 482:32]
  wire  _GEN_403 = invtags_1 != vtag_15 | _GEN_402; // @[Sbuffer.scala 486:42 493:34]
  wire  _sameBlockInflightMask_mask_T_33 = stateVec_0_state_inflight & _T_86; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_35 = stateVec_1_state_inflight & _T_88; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_37 = stateVec_2_state_inflight & _T_90; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_39 = stateVec_3_state_inflight & _T_92; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_41 = stateVec_4_state_inflight & _T_94; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_43 = stateVec_5_state_inflight & _T_96; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_45 = stateVec_6_state_inflight & _T_98; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_47 = stateVec_7_state_inflight & _T_100; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_49 = stateVec_8_state_inflight & _T_102; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_51 = stateVec_9_state_inflight & _T_104; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_53 = stateVec_10_state_inflight & _T_106; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_55 = stateVec_11_state_inflight & _T_108; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_57 = stateVec_12_state_inflight & _T_110; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_59 = stateVec_13_state_inflight & _T_112; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_61 = stateVec_14_state_inflight & _T_114; // @[Sbuffer.scala 599:54]
  wire  _sameBlockInflightMask_mask_T_63 = stateVec_15_state_inflight & _T_116; // @[Sbuffer.scala 599:54]
  wire [7:0] sameBlockInflightMask_mask_lo_1 = {_sameBlockInflightMask_mask_T_47,_sameBlockInflightMask_mask_T_45,
    _sameBlockInflightMask_mask_T_43,_sameBlockInflightMask_mask_T_41,_sameBlockInflightMask_mask_T_39,
    _sameBlockInflightMask_mask_T_37,_sameBlockInflightMask_mask_T_35,_sameBlockInflightMask_mask_T_33}; // @[Sbuffer.scala 599:79]
  wire [15:0] sameBlockInflightMask_1 = {_sameBlockInflightMask_mask_T_63,_sameBlockInflightMask_mask_T_61,
    _sameBlockInflightMask_mask_T_59,_sameBlockInflightMask_mask_T_57,_sameBlockInflightMask_mask_T_55,
    _sameBlockInflightMask_mask_T_53,_sameBlockInflightMask_mask_T_51,_sameBlockInflightMask_mask_T_49,
    sameBlockInflightMask_mask_lo_1}; // @[Sbuffer.scala 599:79]
  wire  _stateVec_0_w_sameblock_inflight_T_1 = |sameBlockInflightMask_1; // @[Sbuffer.scala 460:74]
  wire  _GEN_407 = secondInsertVec[0] | _GEN_278; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_408 = secondInsertVec[0] ? |sameBlockInflightMask_1 : _GEN_279; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_414 = secondInsertVec[1] | _GEN_283; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_415 = secondInsertVec[1] ? |sameBlockInflightMask_1 : _GEN_284; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_421 = secondInsertVec[2] | _GEN_288; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_422 = secondInsertVec[2] ? |sameBlockInflightMask_1 : _GEN_289; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_428 = secondInsertVec[3] | _GEN_293; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_429 = secondInsertVec[3] ? |sameBlockInflightMask_1 : _GEN_294; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_435 = secondInsertVec[4] | _GEN_298; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_436 = secondInsertVec[4] ? |sameBlockInflightMask_1 : _GEN_299; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_442 = secondInsertVec[5] | _GEN_303; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_443 = secondInsertVec[5] ? |sameBlockInflightMask_1 : _GEN_304; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_449 = secondInsertVec[6] | _GEN_308; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_450 = secondInsertVec[6] ? |sameBlockInflightMask_1 : _GEN_309; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_456 = secondInsertVec[7] | _GEN_313; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_457 = secondInsertVec[7] ? |sameBlockInflightMask_1 : _GEN_314; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_463 = secondInsertVec[8] | _GEN_318; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_464 = secondInsertVec[8] ? |sameBlockInflightMask_1 : _GEN_319; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_470 = secondInsertVec[9] | _GEN_323; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_471 = secondInsertVec[9] ? |sameBlockInflightMask_1 : _GEN_324; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_477 = secondInsertVec[10] | _GEN_328; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_478 = secondInsertVec[10] ? |sameBlockInflightMask_1 : _GEN_329; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_484 = secondInsertVec[11] | _GEN_333; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_485 = secondInsertVec[11] ? |sameBlockInflightMask_1 : _GEN_334; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_491 = secondInsertVec[12] | _GEN_338; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_492 = secondInsertVec[12] ? |sameBlockInflightMask_1 : _GEN_339; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_498 = secondInsertVec[13] | _GEN_343; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_499 = secondInsertVec[13] ? |sameBlockInflightMask_1 : _GEN_344; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_505 = secondInsertVec[14] | _GEN_348; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_506 = secondInsertVec[14] ? |sameBlockInflightMask_1 : _GEN_349; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_512 = secondInsertVec[15] | _GEN_353; // @[Sbuffer.scala 458:32 459:40]
  wire  _GEN_513 = secondInsertVec[15] ? |sameBlockInflightMask_1 : _GEN_354; // @[Sbuffer.scala 458:32 460:49]
  wire  _GEN_536 = canMerge_1 ? _GEN_278 : _GEN_407; // @[Sbuffer.scala 512:24]
  wire  _GEN_541 = canMerge_1 ? _GEN_283 : _GEN_414; // @[Sbuffer.scala 512:24]
  wire  _GEN_546 = canMerge_1 ? _GEN_288 : _GEN_421; // @[Sbuffer.scala 512:24]
  wire  _GEN_551 = canMerge_1 ? _GEN_293 : _GEN_428; // @[Sbuffer.scala 512:24]
  wire  _GEN_556 = canMerge_1 ? _GEN_298 : _GEN_435; // @[Sbuffer.scala 512:24]
  wire  _GEN_561 = canMerge_1 ? _GEN_303 : _GEN_442; // @[Sbuffer.scala 512:24]
  wire  _GEN_566 = canMerge_1 ? _GEN_308 : _GEN_449; // @[Sbuffer.scala 512:24]
  wire  _GEN_571 = canMerge_1 ? _GEN_313 : _GEN_456; // @[Sbuffer.scala 512:24]
  wire  _GEN_576 = canMerge_1 ? _GEN_318 : _GEN_463; // @[Sbuffer.scala 512:24]
  wire  _GEN_581 = canMerge_1 ? _GEN_323 : _GEN_470; // @[Sbuffer.scala 512:24]
  wire  _GEN_586 = canMerge_1 ? _GEN_328 : _GEN_477; // @[Sbuffer.scala 512:24]
  wire  _GEN_591 = canMerge_1 ? _GEN_333 : _GEN_484; // @[Sbuffer.scala 512:24]
  wire  _GEN_596 = canMerge_1 ? _GEN_338 : _GEN_491; // @[Sbuffer.scala 512:24]
  wire  _GEN_601 = canMerge_1 ? _GEN_343 : _GEN_498; // @[Sbuffer.scala 512:24]
  wire  _GEN_606 = canMerge_1 ? _GEN_348 : _GEN_505; // @[Sbuffer.scala 512:24]
  wire  _GEN_611 = canMerge_1 ? _GEN_353 : _GEN_512; // @[Sbuffer.scala 512:24]
  wire  _GEN_634 = _dataModule_io_writeReq_1_valid_T ? _GEN_536 : _GEN_278; // @[Sbuffer.scala 511:20]
  wire  _GEN_639 = _dataModule_io_writeReq_1_valid_T ? _GEN_541 : _GEN_283; // @[Sbuffer.scala 511:20]
  wire  _GEN_644 = _dataModule_io_writeReq_1_valid_T ? _GEN_546 : _GEN_288; // @[Sbuffer.scala 511:20]
  wire  _GEN_649 = _dataModule_io_writeReq_1_valid_T ? _GEN_551 : _GEN_293; // @[Sbuffer.scala 511:20]
  wire  _GEN_654 = _dataModule_io_writeReq_1_valid_T ? _GEN_556 : _GEN_298; // @[Sbuffer.scala 511:20]
  wire  _GEN_659 = _dataModule_io_writeReq_1_valid_T ? _GEN_561 : _GEN_303; // @[Sbuffer.scala 511:20]
  wire  _GEN_664 = _dataModule_io_writeReq_1_valid_T ? _GEN_566 : _GEN_308; // @[Sbuffer.scala 511:20]
  wire  _GEN_669 = _dataModule_io_writeReq_1_valid_T ? _GEN_571 : _GEN_313; // @[Sbuffer.scala 511:20]
  wire  _GEN_674 = _dataModule_io_writeReq_1_valid_T ? _GEN_576 : _GEN_318; // @[Sbuffer.scala 511:20]
  wire  _GEN_679 = _dataModule_io_writeReq_1_valid_T ? _GEN_581 : _GEN_323; // @[Sbuffer.scala 511:20]
  wire  _GEN_684 = _dataModule_io_writeReq_1_valid_T ? _GEN_586 : _GEN_328; // @[Sbuffer.scala 511:20]
  wire  _GEN_689 = _dataModule_io_writeReq_1_valid_T ? _GEN_591 : _GEN_333; // @[Sbuffer.scala 511:20]
  wire  _GEN_694 = _dataModule_io_writeReq_1_valid_T ? _GEN_596 : _GEN_338; // @[Sbuffer.scala 511:20]
  wire  _GEN_699 = _dataModule_io_writeReq_1_valid_T ? _GEN_601 : _GEN_343; // @[Sbuffer.scala 511:20]
  wire  _GEN_704 = _dataModule_io_writeReq_1_valid_T ? _GEN_606 : _GEN_348; // @[Sbuffer.scala 511:20]
  wire  _GEN_709 = _dataModule_io_writeReq_1_valid_T ? _GEN_611 : _GEN_353; // @[Sbuffer.scala 511:20]
  wire [7:0] sbuffer_empty_lo = {invalidMask_8,invalidMask_9,invalidMask_10,invalidMask_11,invalidMask_12,invalidMask_13
    ,invalidMask_14,invalidMask_15}; // @[Cat.scala 33:92]
  wire [15:0] _sbuffer_empty_T = {invalidMask_0,invalidMask_1,invalidMask_2,invalidMask_3,invalidMask_4,invalidMask_5,
    invalidMask_6,invalidMask_7,sbuffer_empty_lo}; // @[Cat.scala 33:92]
  wire  sbuffer_empty = &_sbuffer_empty_T; // @[Sbuffer.scala 546:44]
  wire [1:0] _sq_empty_T = {io_in_0_valid,io_in_1_valid}; // @[Cat.scala 33:92]
  wire  sq_empty = ~(|_sq_empty_T); // @[Sbuffer.scala 547:18]
  wire  empty = sbuffer_empty & sq_empty; // @[Sbuffer.scala 548:29]
  reg [4:0] threshold; // @[Sbuffer.scala 549:26]
  wire [1:0] _ActiveCount_T = _candidateVec_T_1 + _candidateVec_T_5; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_2 = _candidateVec_T_9 + _candidateVec_T_13; // @[Bitwise.scala 51:90]
  wire [2:0] _ActiveCount_T_4 = _ActiveCount_T + _ActiveCount_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_6 = _candidateVec_T_17 + _candidateVec_T_21; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_8 = _candidateVec_T_25 + _candidateVec_T_29; // @[Bitwise.scala 51:90]
  wire [2:0] _ActiveCount_T_10 = _ActiveCount_T_6 + _ActiveCount_T_8; // @[Bitwise.scala 51:90]
  wire [3:0] _ActiveCount_T_12 = _ActiveCount_T_4 + _ActiveCount_T_10; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_14 = _candidateVec_T_33 + _candidateVec_T_37; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_16 = _candidateVec_T_41 + _candidateVec_T_45; // @[Bitwise.scala 51:90]
  wire [2:0] _ActiveCount_T_18 = _ActiveCount_T_14 + _ActiveCount_T_16; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_20 = _candidateVec_T_49 + _candidateVec_T_53; // @[Bitwise.scala 51:90]
  wire [1:0] _ActiveCount_T_22 = _candidateVec_T_57 + _candidateVec_T_61; // @[Bitwise.scala 51:90]
  wire [2:0] _ActiveCount_T_24 = _ActiveCount_T_20 + _ActiveCount_T_22; // @[Bitwise.scala 51:90]
  wire [3:0] _ActiveCount_T_26 = _ActiveCount_T_18 + _ActiveCount_T_24; // @[Bitwise.scala 51:90]
  wire [4:0] ActiveCount = _ActiveCount_T_12 + _ActiveCount_T_26; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T = stateVec_0_state_valid + stateVec_1_state_valid; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_2 = stateVec_2_state_valid + stateVec_3_state_valid; // @[Bitwise.scala 51:90]
  wire [2:0] _ValidCount_T_4 = _ValidCount_T + _ValidCount_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_6 = stateVec_4_state_valid + stateVec_5_state_valid; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_8 = stateVec_6_state_valid + stateVec_7_state_valid; // @[Bitwise.scala 51:90]
  wire [2:0] _ValidCount_T_10 = _ValidCount_T_6 + _ValidCount_T_8; // @[Bitwise.scala 51:90]
  wire [3:0] _ValidCount_T_12 = _ValidCount_T_4 + _ValidCount_T_10; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_14 = stateVec_8_state_valid + stateVec_9_state_valid; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_16 = stateVec_10_state_valid + stateVec_11_state_valid; // @[Bitwise.scala 51:90]
  wire [2:0] _ValidCount_T_18 = _ValidCount_T_14 + _ValidCount_T_16; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_20 = stateVec_12_state_valid + stateVec_13_state_valid; // @[Bitwise.scala 51:90]
  wire [1:0] _ValidCount_T_22 = stateVec_14_state_valid + stateVec_15_state_valid; // @[Bitwise.scala 51:90]
  wire [2:0] _ValidCount_T_24 = _ValidCount_T_20 + _ValidCount_T_22; // @[Bitwise.scala 51:90]
  wire [3:0] _ValidCount_T_26 = _ValidCount_T_18 + _ValidCount_T_24; // @[Bitwise.scala 51:90]
  wire [4:0] ValidCount = _ValidCount_T_12 + _ValidCount_T_26; // @[Bitwise.scala 51:90]
  reg  do_eviction; // @[Sbuffer.scala 552:28]
  reg  io_flush_empty_REG; // @[Sbuffer.scala 557:28]
  wire [1:0] _GEN_718 = sbuffer_empty ? 2'h0 : sbuffer_state; // @[Sbuffer.scala 577:32 578:23 295:30]
  wire [1:0] _GEN_720 = ~do_eviction ? 2'h0 : sbuffer_state; // @[Sbuffer.scala 586:31 587:23 295:30]
  wire [1:0] _GEN_721 = do_uarch_drain ? 2'h3 : _GEN_720; // @[Sbuffer.scala 584:33 585:23]
  wire [1:0] _GEN_722 = io_flush_valid ? 2'h2 : _GEN_721; // @[Sbuffer.scala 582:27 583:23]
  wire  need_drain = sbuffer_state[1]; // @[Sbuffer.scala 294:10]
  wire  need_replace = do_eviction | sbuffer_state == 2'h1; // @[Sbuffer.scala 633:34]
  wire [3:0] _sbuffer_out_s0_evictionIdx_T = cohHasTimeOut ? cohTimeOutIdx : Sbuffer_PLRU_io_replaceWay; // @[Sbuffer.scala 638:10]
  wire [3:0] _sbuffer_out_s0_evictionIdx_T_1 = need_drain ? drainIdx : _sbuffer_out_s0_evictionIdx_T; // @[Sbuffer.scala 636:8]
  wire [3:0] sbuffer_out_s0_evictionIdx = missqReplayHasTimeOut ? missqReplayTimeOutIdx :
    _sbuffer_out_s0_evictionIdx_T_1; // @[Sbuffer.scala 634:39]
  wire  _GEN_728 = 4'h1 == sbuffer_out_s0_evictionIdx ? stateVec_1_state_inflight : stateVec_0_state_inflight; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_729 = 4'h2 == sbuffer_out_s0_evictionIdx ? stateVec_2_state_inflight : _GEN_728; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_730 = 4'h3 == sbuffer_out_s0_evictionIdx ? stateVec_3_state_inflight : _GEN_729; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_731 = 4'h4 == sbuffer_out_s0_evictionIdx ? stateVec_4_state_inflight : _GEN_730; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_732 = 4'h5 == sbuffer_out_s0_evictionIdx ? stateVec_5_state_inflight : _GEN_731; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_733 = 4'h6 == sbuffer_out_s0_evictionIdx ? stateVec_6_state_inflight : _GEN_732; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_734 = 4'h7 == sbuffer_out_s0_evictionIdx ? stateVec_7_state_inflight : _GEN_733; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_735 = 4'h8 == sbuffer_out_s0_evictionIdx ? stateVec_8_state_inflight : _GEN_734; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_736 = 4'h9 == sbuffer_out_s0_evictionIdx ? stateVec_9_state_inflight : _GEN_735; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_737 = 4'ha == sbuffer_out_s0_evictionIdx ? stateVec_10_state_inflight : _GEN_736; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_738 = 4'hb == sbuffer_out_s0_evictionIdx ? stateVec_11_state_inflight : _GEN_737; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_739 = 4'hc == sbuffer_out_s0_evictionIdx ? stateVec_12_state_inflight : _GEN_738; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_740 = 4'hd == sbuffer_out_s0_evictionIdx ? stateVec_13_state_inflight : _GEN_739; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_741 = 4'he == sbuffer_out_s0_evictionIdx ? stateVec_14_state_inflight : _GEN_740; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_742 = 4'hf == sbuffer_out_s0_evictionIdx ? stateVec_15_state_inflight : _GEN_741; // @[Sbuffer.scala 66:{53,53}]
  wire  _GEN_744 = 4'h1 == sbuffer_out_s0_evictionIdx ? stateVec_1_state_valid : stateVec_0_state_valid; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_745 = 4'h2 == sbuffer_out_s0_evictionIdx ? stateVec_2_state_valid : _GEN_744; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_746 = 4'h3 == sbuffer_out_s0_evictionIdx ? stateVec_3_state_valid : _GEN_745; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_747 = 4'h4 == sbuffer_out_s0_evictionIdx ? stateVec_4_state_valid : _GEN_746; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_748 = 4'h5 == sbuffer_out_s0_evictionIdx ? stateVec_5_state_valid : _GEN_747; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_749 = 4'h6 == sbuffer_out_s0_evictionIdx ? stateVec_6_state_valid : _GEN_748; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_750 = 4'h7 == sbuffer_out_s0_evictionIdx ? stateVec_7_state_valid : _GEN_749; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_751 = 4'h8 == sbuffer_out_s0_evictionIdx ? stateVec_8_state_valid : _GEN_750; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_752 = 4'h9 == sbuffer_out_s0_evictionIdx ? stateVec_9_state_valid : _GEN_751; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_753 = 4'ha == sbuffer_out_s0_evictionIdx ? stateVec_10_state_valid : _GEN_752; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_754 = 4'hb == sbuffer_out_s0_evictionIdx ? stateVec_11_state_valid : _GEN_753; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_755 = 4'hc == sbuffer_out_s0_evictionIdx ? stateVec_12_state_valid : _GEN_754; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_756 = 4'hd == sbuffer_out_s0_evictionIdx ? stateVec_13_state_valid : _GEN_755; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_757 = 4'he == sbuffer_out_s0_evictionIdx ? stateVec_14_state_valid : _GEN_756; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_758 = 4'hf == sbuffer_out_s0_evictionIdx ? stateVec_15_state_valid : _GEN_757; // @[Sbuffer.scala 66:{50,50}]
  wire  _GEN_760 = 4'h1 == sbuffer_out_s0_evictionIdx ? stateVec_1_w_sameblock_inflight :
    stateVec_0_w_sameblock_inflight; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_761 = 4'h2 == sbuffer_out_s0_evictionIdx ? stateVec_2_w_sameblock_inflight : _GEN_760; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_762 = 4'h3 == sbuffer_out_s0_evictionIdx ? stateVec_3_w_sameblock_inflight : _GEN_761; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_763 = 4'h4 == sbuffer_out_s0_evictionIdx ? stateVec_4_w_sameblock_inflight : _GEN_762; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_764 = 4'h5 == sbuffer_out_s0_evictionIdx ? stateVec_5_w_sameblock_inflight : _GEN_763; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_765 = 4'h6 == sbuffer_out_s0_evictionIdx ? stateVec_6_w_sameblock_inflight : _GEN_764; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_766 = 4'h7 == sbuffer_out_s0_evictionIdx ? stateVec_7_w_sameblock_inflight : _GEN_765; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_767 = 4'h8 == sbuffer_out_s0_evictionIdx ? stateVec_8_w_sameblock_inflight : _GEN_766; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_768 = 4'h9 == sbuffer_out_s0_evictionIdx ? stateVec_9_w_sameblock_inflight : _GEN_767; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_769 = 4'ha == sbuffer_out_s0_evictionIdx ? stateVec_10_w_sameblock_inflight : _GEN_768; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_770 = 4'hb == sbuffer_out_s0_evictionIdx ? stateVec_11_w_sameblock_inflight : _GEN_769; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_771 = 4'hc == sbuffer_out_s0_evictionIdx ? stateVec_12_w_sameblock_inflight : _GEN_770; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_772 = 4'hd == sbuffer_out_s0_evictionIdx ? stateVec_13_w_sameblock_inflight : _GEN_771; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_773 = 4'he == sbuffer_out_s0_evictionIdx ? stateVec_14_w_sameblock_inflight : _GEN_772; // @[Sbuffer.scala 66:{72,72}]
  wire  _GEN_774 = 4'hf == sbuffer_out_s0_evictionIdx ? stateVec_15_w_sameblock_inflight : _GEN_773; // @[Sbuffer.scala 66:{72,72}]
  wire  _sbuffer_out_s0_valid_T_3 = _GEN_758 & ~_GEN_742 & ~_GEN_774; // @[Sbuffer.scala 66:69]
  wire  _sbuffer_out_s0_valid_T_5 = need_drain | cohHasTimeOut | need_replace; // @[Sbuffer.scala 646:34]
  wire  _sbuffer_out_s0_valid_T_6 = _sbuffer_out_s0_valid_T_3 & _sbuffer_out_s0_valid_T_5; // @[Sbuffer.scala 645:65]
  wire  sbuffer_out_s0_valid = missqReplayHasTimeOut | _sbuffer_out_s0_valid_T_6; // @[Sbuffer.scala 644:52]
  wire [29:0] _GEN_776 = 4'h1 == sbuffer_out_s0_evictionIdx ? ptag_1 : ptag_0; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_777 = 4'h2 == sbuffer_out_s0_evictionIdx ? ptag_2 : _GEN_776; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_778 = 4'h3 == sbuffer_out_s0_evictionIdx ? ptag_3 : _GEN_777; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_779 = 4'h4 == sbuffer_out_s0_evictionIdx ? ptag_4 : _GEN_778; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_780 = 4'h5 == sbuffer_out_s0_evictionIdx ? ptag_5 : _GEN_779; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_781 = 4'h6 == sbuffer_out_s0_evictionIdx ? ptag_6 : _GEN_780; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_782 = 4'h7 == sbuffer_out_s0_evictionIdx ? ptag_7 : _GEN_781; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_783 = 4'h8 == sbuffer_out_s0_evictionIdx ? ptag_8 : _GEN_782; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_784 = 4'h9 == sbuffer_out_s0_evictionIdx ? ptag_9 : _GEN_783; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_785 = 4'ha == sbuffer_out_s0_evictionIdx ? ptag_10 : _GEN_784; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_786 = 4'hb == sbuffer_out_s0_evictionIdx ? ptag_11 : _GEN_785; // @[Sbuffer.scala 595:{53,53}]
  wire [29:0] _GEN_787 = 4'hc == sbuffer_out_s0_evictionIdx ? ptag_12 : _GEN_786; // @[Sbuffer.scala 595:{53,53}]
  reg  blockDcacheWrite; // @[Sbuffer.scala 659:38]
  wire  _sbuffer_out_s1_ready_T = ~blockDcacheWrite; // @[Sbuffer.scala 667:50]
  reg  sbuffer_out_s1_valid; // @[Sbuffer.scala 666:37]
  wire  sbuffer_out_s0_cango = io_dcache_req_ready & ~blockDcacheWrite | ~sbuffer_out_s1_valid; // @[Sbuffer.scala 667:68]
  wire  sbuffer_out_s0_fire = sbuffer_out_s0_valid & sbuffer_out_s0_cango; // @[Sbuffer.scala 652:47]
  wire [15:0] _shouldWaitWriteFinish_T = 16'h1 << sbuffer_out_s0_evictionIdx; // @[OneHot.scala 57:35]
  wire [15:0] _shouldWaitWriteFinish_T_1 = dataModule_io_writeReq_0_bits_wvec & _shouldWaitWriteFinish_T; // @[Sbuffer.scala 660:35]
  wire  _shouldWaitWriteFinish_T_3 = |_shouldWaitWriteFinish_T_1 & dataModule_io_writeReq_0_valid; // @[Sbuffer.scala 660:86]
  wire [15:0] _shouldWaitWriteFinish_T_5 = dataModule_io_writeReq_1_bits_wvec & _shouldWaitWriteFinish_T; // @[Sbuffer.scala 660:35]
  wire  _shouldWaitWriteFinish_T_7 = |_shouldWaitWriteFinish_T_5 & dataModule_io_writeReq_1_valid; // @[Sbuffer.scala 660:86]
  wire [1:0] _shouldWaitWriteFinish_T_8 = {_shouldWaitWriteFinish_T_7,_shouldWaitWriteFinish_T_3}; // @[Sbuffer.scala 662:6]
  wire  sbuffer_out_s1_fire = io_dcache_req_ready & io_dcache_req_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_793 = 4'h0 == sbuffer_out_s0_evictionIdx | stateVec_0_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_794 = 4'h1 == sbuffer_out_s0_evictionIdx | stateVec_1_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_795 = 4'h2 == sbuffer_out_s0_evictionIdx | stateVec_2_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_796 = 4'h3 == sbuffer_out_s0_evictionIdx | stateVec_3_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_797 = 4'h4 == sbuffer_out_s0_evictionIdx | stateVec_4_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_798 = 4'h5 == sbuffer_out_s0_evictionIdx | stateVec_5_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_799 = 4'h6 == sbuffer_out_s0_evictionIdx | stateVec_6_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_800 = 4'h7 == sbuffer_out_s0_evictionIdx | stateVec_7_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_801 = 4'h8 == sbuffer_out_s0_evictionIdx | stateVec_8_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_802 = 4'h9 == sbuffer_out_s0_evictionIdx | stateVec_9_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_803 = 4'ha == sbuffer_out_s0_evictionIdx | stateVec_10_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_804 = 4'hb == sbuffer_out_s0_evictionIdx | stateVec_11_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_805 = 4'hc == sbuffer_out_s0_evictionIdx | stateVec_12_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_806 = 4'hd == sbuffer_out_s0_evictionIdx | stateVec_13_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_807 = 4'he == sbuffer_out_s0_evictionIdx | stateVec_14_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_808 = 4'hf == sbuffer_out_s0_evictionIdx | stateVec_15_state_inflight; // @[Sbuffer.scala 280:25 679:{57,57}]
  wire  _GEN_809 = 4'h0 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_0_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_810 = 4'h1 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_1_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_811 = 4'h2 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_2_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_812 = 4'h3 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_3_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_813 = 4'h4 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_4_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_814 = 4'h5 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_5_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_815 = 4'h6 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_6_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_816 = 4'h7 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_7_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_817 = 4'h8 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_8_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_818 = 4'h9 == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_9_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_819 = 4'ha == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_10_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_820 = 4'hb == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_11_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_821 = 4'hc == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_12_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_822 = 4'hd == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_13_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_823 = 4'he == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_14_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_824 = 4'hf == sbuffer_out_s0_evictionIdx ? 1'h0 : stateVec_15_w_timeout; // @[Sbuffer.scala 280:25 680:{52,52}]
  wire  _GEN_825 = sbuffer_out_s0_fire ? _GEN_793 : stateVec_0_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_826 = sbuffer_out_s0_fire ? _GEN_794 : stateVec_1_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_827 = sbuffer_out_s0_fire ? _GEN_795 : stateVec_2_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_828 = sbuffer_out_s0_fire ? _GEN_796 : stateVec_3_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_829 = sbuffer_out_s0_fire ? _GEN_797 : stateVec_4_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_830 = sbuffer_out_s0_fire ? _GEN_798 : stateVec_5_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_831 = sbuffer_out_s0_fire ? _GEN_799 : stateVec_6_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_832 = sbuffer_out_s0_fire ? _GEN_800 : stateVec_7_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_833 = sbuffer_out_s0_fire ? _GEN_801 : stateVec_8_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_834 = sbuffer_out_s0_fire ? _GEN_802 : stateVec_9_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_835 = sbuffer_out_s0_fire ? _GEN_803 : stateVec_10_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_836 = sbuffer_out_s0_fire ? _GEN_804 : stateVec_11_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_837 = sbuffer_out_s0_fire ? _GEN_805 : stateVec_12_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_838 = sbuffer_out_s0_fire ? _GEN_806 : stateVec_13_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_839 = sbuffer_out_s0_fire ? _GEN_807 : stateVec_14_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_840 = sbuffer_out_s0_fire ? _GEN_808 : stateVec_15_state_inflight; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_841 = sbuffer_out_s0_fire ? _GEN_809 : stateVec_0_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_842 = sbuffer_out_s0_fire ? _GEN_810 : stateVec_1_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_843 = sbuffer_out_s0_fire ? _GEN_811 : stateVec_2_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_844 = sbuffer_out_s0_fire ? _GEN_812 : stateVec_3_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_845 = sbuffer_out_s0_fire ? _GEN_813 : stateVec_4_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_846 = sbuffer_out_s0_fire ? _GEN_814 : stateVec_5_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_847 = sbuffer_out_s0_fire ? _GEN_815 : stateVec_6_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_848 = sbuffer_out_s0_fire ? _GEN_816 : stateVec_7_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_849 = sbuffer_out_s0_fire ? _GEN_817 : stateVec_8_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_850 = sbuffer_out_s0_fire ? _GEN_818 : stateVec_9_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_851 = sbuffer_out_s0_fire ? _GEN_819 : stateVec_10_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_852 = sbuffer_out_s0_fire ? _GEN_820 : stateVec_11_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_853 = sbuffer_out_s0_fire ? _GEN_821 : stateVec_12_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_854 = sbuffer_out_s0_fire ? _GEN_822 : stateVec_13_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_855 = sbuffer_out_s0_fire ? _GEN_823 : stateVec_14_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_856 = sbuffer_out_s0_fire ? _GEN_824 : stateVec_15_w_timeout; // @[Sbuffer.scala 280:25 678:28]
  wire  _GEN_858 = 4'h1 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_5 : _candidateVec_T_1; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_859 = 4'h2 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_9 : _GEN_858; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_860 = 4'h3 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_13 : _GEN_859; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_861 = 4'h4 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_17 : _GEN_860; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_862 = 4'h5 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_21 : _GEN_861; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_863 = 4'h6 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_25 : _GEN_862; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_864 = 4'h7 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_29 : _GEN_863; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_865 = 4'h8 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_33 : _GEN_864; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_866 = 4'h9 == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_37 : _GEN_865; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_867 = 4'ha == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_41 : _GEN_866; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_868 = 4'hb == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_45 : _GEN_867; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_869 = 4'hc == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_49 : _GEN_868; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_870 = 4'hd == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_53 : _GEN_869; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_871 = 4'he == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_57 : _GEN_870; // @[Sbuffer.scala 692:{101,101}]
  wire  _GEN_872 = 4'hf == Sbuffer_PLRU_io_replaceWay ? _candidateVec_T_61 : _GEN_871; // @[Sbuffer.scala 692:{101,101}]
  wire  _accessIdx_2_valid_T_7 = need_replace & ~need_drain & ~cohHasTimeOut & ~missqReplayHasTimeOut &
    sbuffer_out_s0_cango & _GEN_872; // @[Sbuffer.scala 692:101]
  wire  _GEN_874 = 4'h1 == Sbuffer_PLRU_io_replaceWay ? invalidMask_1 : invalidMask_0; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_875 = 4'h2 == Sbuffer_PLRU_io_replaceWay ? invalidMask_2 : _GEN_874; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_876 = 4'h3 == Sbuffer_PLRU_io_replaceWay ? invalidMask_3 : _GEN_875; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_877 = 4'h4 == Sbuffer_PLRU_io_replaceWay ? invalidMask_4 : _GEN_876; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_878 = 4'h5 == Sbuffer_PLRU_io_replaceWay ? invalidMask_5 : _GEN_877; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_879 = 4'h6 == Sbuffer_PLRU_io_replaceWay ? invalidMask_6 : _GEN_878; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_880 = 4'h7 == Sbuffer_PLRU_io_replaceWay ? invalidMask_7 : _GEN_879; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_881 = 4'h8 == Sbuffer_PLRU_io_replaceWay ? invalidMask_8 : _GEN_880; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_882 = 4'h9 == Sbuffer_PLRU_io_replaceWay ? invalidMask_9 : _GEN_881; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_883 = 4'ha == Sbuffer_PLRU_io_replaceWay ? invalidMask_10 : _GEN_882; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_884 = 4'hb == Sbuffer_PLRU_io_replaceWay ? invalidMask_11 : _GEN_883; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_885 = 4'hc == Sbuffer_PLRU_io_replaceWay ? invalidMask_12 : _GEN_884; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_886 = 4'hd == Sbuffer_PLRU_io_replaceWay ? invalidMask_13 : _GEN_885; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_887 = 4'he == Sbuffer_PLRU_io_replaceWay ? invalidMask_14 : _GEN_886; // @[Sbuffer.scala 691:{62,62}]
  wire  _GEN_888 = 4'hf == Sbuffer_PLRU_io_replaceWay ? invalidMask_15 : _GEN_887; // @[Sbuffer.scala 691:{62,62}]
  reg [3:0] sbuffer_out_s1_evictionIdx; // @[Reg.scala 19:16]
  reg [29:0] sbuffer_out_s1_evictionPTag; // @[Reg.scala 19:16]
  reg [32:0] sbuffer_out_s1_evictionVTag; // @[Reg.scala 19:16]
  wire [32:0] _GEN_892 = 4'h1 == sbuffer_out_s0_evictionIdx ? vtag_1 : vtag_0; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_893 = 4'h2 == sbuffer_out_s0_evictionIdx ? vtag_2 : _GEN_892; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_894 = 4'h3 == sbuffer_out_s0_evictionIdx ? vtag_3 : _GEN_893; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_895 = 4'h4 == sbuffer_out_s0_evictionIdx ? vtag_4 : _GEN_894; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_896 = 4'h5 == sbuffer_out_s0_evictionIdx ? vtag_5 : _GEN_895; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_897 = 4'h6 == sbuffer_out_s0_evictionIdx ? vtag_6 : _GEN_896; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_898 = 4'h7 == sbuffer_out_s0_evictionIdx ? vtag_7 : _GEN_897; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_899 = 4'h8 == sbuffer_out_s0_evictionIdx ? vtag_8 : _GEN_898; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_900 = 4'h9 == sbuffer_out_s0_evictionIdx ? vtag_9 : _GEN_899; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_901 = 4'ha == sbuffer_out_s0_evictionIdx ? vtag_10 : _GEN_900; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_902 = 4'hb == sbuffer_out_s0_evictionIdx ? vtag_11 : _GEN_901; // @[Reg.scala 20:{22,22}]
  wire [32:0] _GEN_903 = 4'hc == sbuffer_out_s0_evictionIdx ? vtag_12 : _GEN_902; // @[Reg.scala 20:{22,22}]
  wire [7:0] _GEN_908 = dataModule_io_dataOut_0_0_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_909 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_1 : _GEN_908; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_910 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_1 : _GEN_909; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_911 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_1 : _GEN_910; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_912 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_1 : _GEN_911; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_913 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_1 : _GEN_912; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_914 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_1 : _GEN_913; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_915 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_1 : _GEN_914; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_916 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_1 : _GEN_915; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_917 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_1 : _GEN_916; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_918 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_1 : _GEN_917; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_919 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_1 : _GEN_918; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_920 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_1 : _GEN_919; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_921 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_1 : _GEN_920; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_922 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_1 : _GEN_921; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_923 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_1 : _GEN_922; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_924 = dataModule_io_dataOut_0_0_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_925 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_0 : _GEN_924; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_926 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_0 : _GEN_925; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_927 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_0 : _GEN_926; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_928 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_0 : _GEN_927; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_929 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_0 : _GEN_928; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_930 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_0 : _GEN_929; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_931 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_0 : _GEN_930; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_932 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_0 : _GEN_931; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_933 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_0 : _GEN_932; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_934 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_0 : _GEN_933; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_935 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_0 : _GEN_934; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_936 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_0 : _GEN_935; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_937 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_0 : _GEN_936; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_938 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_0 : _GEN_937; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_939 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_0 : _GEN_938; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_940 = dataModule_io_dataOut_0_0_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_941 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_3 : _GEN_940; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_942 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_3 : _GEN_941; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_943 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_3 : _GEN_942; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_944 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_3 : _GEN_943; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_945 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_3 : _GEN_944; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_946 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_3 : _GEN_945; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_947 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_3 : _GEN_946; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_948 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_3 : _GEN_947; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_949 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_3 : _GEN_948; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_950 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_3 : _GEN_949; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_951 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_3 : _GEN_950; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_952 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_3 : _GEN_951; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_953 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_3 : _GEN_952; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_954 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_3 : _GEN_953; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_955 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_3 : _GEN_954; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_956 = dataModule_io_dataOut_0_0_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_957 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_2 : _GEN_956; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_958 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_2 : _GEN_957; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_959 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_2 : _GEN_958; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_960 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_2 : _GEN_959; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_961 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_2 : _GEN_960; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_962 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_2 : _GEN_961; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_963 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_2 : _GEN_962; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_964 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_2 : _GEN_963; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_965 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_2 : _GEN_964; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_966 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_2 : _GEN_965; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_967 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_2 : _GEN_966; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_968 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_2 : _GEN_967; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_969 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_2 : _GEN_968; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_970 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_2 : _GEN_969; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_971 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_2 : _GEN_970; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_972 = dataModule_io_dataOut_0_0_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_973 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_5 : _GEN_972; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_974 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_5 : _GEN_973; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_975 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_5 : _GEN_974; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_976 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_5 : _GEN_975; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_977 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_5 : _GEN_976; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_978 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_5 : _GEN_977; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_979 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_5 : _GEN_978; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_980 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_5 : _GEN_979; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_981 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_5 : _GEN_980; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_982 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_5 : _GEN_981; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_983 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_5 : _GEN_982; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_984 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_5 : _GEN_983; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_985 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_5 : _GEN_984; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_986 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_5 : _GEN_985; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_987 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_5 : _GEN_986; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_988 = dataModule_io_dataOut_0_0_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_989 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_4 : _GEN_988; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_990 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_4 : _GEN_989; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_991 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_4 : _GEN_990; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_992 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_4 : _GEN_991; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_993 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_4 : _GEN_992; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_994 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_4 : _GEN_993; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_995 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_4 : _GEN_994; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_996 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_4 : _GEN_995; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_997 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_4 : _GEN_996; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_998 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_4 : _GEN_997; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_999 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_4 : _GEN_998; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1000 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_4 : _GEN_999; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1001 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_4 : _GEN_1000; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1002 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_4 : _GEN_1001; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1003 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_4 : _GEN_1002; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1004 = dataModule_io_dataOut_0_0_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1005 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_7 : _GEN_1004; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1006 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_7 : _GEN_1005; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1007 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_7 : _GEN_1006; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1008 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_7 : _GEN_1007; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1009 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_7 : _GEN_1008; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1010 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_7 : _GEN_1009; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1011 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_7 : _GEN_1010; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1012 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_7 : _GEN_1011; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1013 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_7 : _GEN_1012; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1014 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_7 : _GEN_1013; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1015 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_7 : _GEN_1014; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1016 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_7 : _GEN_1015; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1017 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_7 : _GEN_1016; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1018 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_7 : _GEN_1017; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1019 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_7 : _GEN_1018; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1020 = dataModule_io_dataOut_0_0_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1021 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_0_6 : _GEN_1020; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1022 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_0_6 : _GEN_1021; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1023 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_0_6 : _GEN_1022; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1024 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_0_6 : _GEN_1023; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1025 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_0_6 : _GEN_1024; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1026 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_0_6 : _GEN_1025; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1027 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_0_6 : _GEN_1026; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1028 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_0_6 : _GEN_1027; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1029 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_0_6 : _GEN_1028; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1030 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_0_6 : _GEN_1029; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1031 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_0_6 : _GEN_1030; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1032 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_0_6 : _GEN_1031; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1033 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_0_6 : _GEN_1032; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1034 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_0_6 : _GEN_1033; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1035 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_0_6 : _GEN_1034; // @[Sbuffer.scala 703:{64,64}]
  wire [63:0] io_dcache_req_bits_data_lo_lo_lo = {_GEN_1019,_GEN_1035,_GEN_987,_GEN_1003,_GEN_955,_GEN_971,_GEN_923,
    _GEN_939}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1036 = dataModule_io_dataOut_0_1_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1037 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_1 : _GEN_1036; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1038 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_1 : _GEN_1037; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1039 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_1 : _GEN_1038; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1040 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_1 : _GEN_1039; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1041 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_1 : _GEN_1040; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1042 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_1 : _GEN_1041; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1043 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_1 : _GEN_1042; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1044 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_1 : _GEN_1043; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1045 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_1 : _GEN_1044; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1046 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_1 : _GEN_1045; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1047 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_1 : _GEN_1046; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1048 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_1 : _GEN_1047; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1049 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_1 : _GEN_1048; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1050 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_1 : _GEN_1049; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1051 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_1 : _GEN_1050; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1052 = dataModule_io_dataOut_0_1_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1053 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_0 : _GEN_1052; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1054 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_0 : _GEN_1053; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1055 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_0 : _GEN_1054; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1056 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_0 : _GEN_1055; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1057 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_0 : _GEN_1056; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1058 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_0 : _GEN_1057; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1059 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_0 : _GEN_1058; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1060 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_0 : _GEN_1059; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1061 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_0 : _GEN_1060; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1062 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_0 : _GEN_1061; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1063 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_0 : _GEN_1062; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1064 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_0 : _GEN_1063; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1065 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_0 : _GEN_1064; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1066 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_0 : _GEN_1065; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1067 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_0 : _GEN_1066; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1068 = dataModule_io_dataOut_0_1_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1069 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_3 : _GEN_1068; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1070 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_3 : _GEN_1069; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1071 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_3 : _GEN_1070; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1072 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_3 : _GEN_1071; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1073 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_3 : _GEN_1072; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1074 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_3 : _GEN_1073; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1075 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_3 : _GEN_1074; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1076 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_3 : _GEN_1075; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1077 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_3 : _GEN_1076; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1078 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_3 : _GEN_1077; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1079 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_3 : _GEN_1078; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1080 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_3 : _GEN_1079; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1081 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_3 : _GEN_1080; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1082 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_3 : _GEN_1081; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1083 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_3 : _GEN_1082; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1084 = dataModule_io_dataOut_0_1_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1085 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_2 : _GEN_1084; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1086 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_2 : _GEN_1085; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1087 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_2 : _GEN_1086; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1088 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_2 : _GEN_1087; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1089 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_2 : _GEN_1088; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1090 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_2 : _GEN_1089; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1091 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_2 : _GEN_1090; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1092 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_2 : _GEN_1091; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1093 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_2 : _GEN_1092; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1094 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_2 : _GEN_1093; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1095 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_2 : _GEN_1094; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1096 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_2 : _GEN_1095; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1097 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_2 : _GEN_1096; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1098 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_2 : _GEN_1097; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1099 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_2 : _GEN_1098; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1100 = dataModule_io_dataOut_0_1_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1101 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_5 : _GEN_1100; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1102 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_5 : _GEN_1101; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1103 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_5 : _GEN_1102; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1104 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_5 : _GEN_1103; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1105 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_5 : _GEN_1104; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1106 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_5 : _GEN_1105; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1107 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_5 : _GEN_1106; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1108 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_5 : _GEN_1107; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1109 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_5 : _GEN_1108; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1110 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_5 : _GEN_1109; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1111 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_5 : _GEN_1110; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1112 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_5 : _GEN_1111; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1113 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_5 : _GEN_1112; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1114 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_5 : _GEN_1113; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1115 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_5 : _GEN_1114; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1116 = dataModule_io_dataOut_0_1_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1117 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_4 : _GEN_1116; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1118 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_4 : _GEN_1117; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1119 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_4 : _GEN_1118; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1120 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_4 : _GEN_1119; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1121 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_4 : _GEN_1120; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1122 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_4 : _GEN_1121; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1123 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_4 : _GEN_1122; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1124 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_4 : _GEN_1123; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1125 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_4 : _GEN_1124; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1126 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_4 : _GEN_1125; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1127 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_4 : _GEN_1126; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1128 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_4 : _GEN_1127; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1129 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_4 : _GEN_1128; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1130 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_4 : _GEN_1129; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1131 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_4 : _GEN_1130; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1132 = dataModule_io_dataOut_0_1_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1133 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_7 : _GEN_1132; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1134 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_7 : _GEN_1133; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1135 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_7 : _GEN_1134; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1136 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_7 : _GEN_1135; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1137 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_7 : _GEN_1136; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1138 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_7 : _GEN_1137; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1139 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_7 : _GEN_1138; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1140 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_7 : _GEN_1139; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1141 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_7 : _GEN_1140; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1142 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_7 : _GEN_1141; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1143 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_7 : _GEN_1142; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1144 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_7 : _GEN_1143; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1145 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_7 : _GEN_1144; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1146 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_7 : _GEN_1145; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1147 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_7 : _GEN_1146; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1148 = dataModule_io_dataOut_0_1_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1149 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_1_6 : _GEN_1148; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1150 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_1_6 : _GEN_1149; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1151 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_1_6 : _GEN_1150; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1152 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_1_6 : _GEN_1151; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1153 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_1_6 : _GEN_1152; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1154 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_1_6 : _GEN_1153; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1155 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_1_6 : _GEN_1154; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1156 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_1_6 : _GEN_1155; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1157 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_1_6 : _GEN_1156; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1158 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_1_6 : _GEN_1157; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1159 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_1_6 : _GEN_1158; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1160 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_1_6 : _GEN_1159; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1161 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_1_6 : _GEN_1160; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1162 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_1_6 : _GEN_1161; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1163 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_1_6 : _GEN_1162; // @[Sbuffer.scala 703:{64,64}]
  wire [127:0] io_dcache_req_bits_data_lo_lo = {_GEN_1147,_GEN_1163,_GEN_1115,_GEN_1131,_GEN_1083,_GEN_1099,_GEN_1051,
    _GEN_1067,io_dcache_req_bits_data_lo_lo_lo}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1164 = dataModule_io_dataOut_0_2_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1165 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_1 : _GEN_1164; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1166 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_1 : _GEN_1165; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1167 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_1 : _GEN_1166; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1168 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_1 : _GEN_1167; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1169 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_1 : _GEN_1168; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1170 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_1 : _GEN_1169; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1171 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_1 : _GEN_1170; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1172 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_1 : _GEN_1171; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1173 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_1 : _GEN_1172; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1174 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_1 : _GEN_1173; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1175 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_1 : _GEN_1174; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1176 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_1 : _GEN_1175; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1177 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_1 : _GEN_1176; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1178 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_1 : _GEN_1177; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1179 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_1 : _GEN_1178; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1180 = dataModule_io_dataOut_0_2_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1181 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_0 : _GEN_1180; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1182 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_0 : _GEN_1181; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1183 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_0 : _GEN_1182; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1184 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_0 : _GEN_1183; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1185 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_0 : _GEN_1184; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1186 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_0 : _GEN_1185; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1187 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_0 : _GEN_1186; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1188 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_0 : _GEN_1187; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1189 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_0 : _GEN_1188; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1190 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_0 : _GEN_1189; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1191 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_0 : _GEN_1190; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1192 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_0 : _GEN_1191; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1193 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_0 : _GEN_1192; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1194 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_0 : _GEN_1193; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1195 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_0 : _GEN_1194; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1196 = dataModule_io_dataOut_0_2_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1197 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_3 : _GEN_1196; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1198 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_3 : _GEN_1197; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1199 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_3 : _GEN_1198; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1200 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_3 : _GEN_1199; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1201 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_3 : _GEN_1200; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1202 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_3 : _GEN_1201; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1203 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_3 : _GEN_1202; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1204 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_3 : _GEN_1203; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1205 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_3 : _GEN_1204; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1206 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_3 : _GEN_1205; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1207 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_3 : _GEN_1206; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1208 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_3 : _GEN_1207; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1209 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_3 : _GEN_1208; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1210 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_3 : _GEN_1209; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1211 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_3 : _GEN_1210; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1212 = dataModule_io_dataOut_0_2_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1213 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_2 : _GEN_1212; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1214 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_2 : _GEN_1213; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1215 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_2 : _GEN_1214; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1216 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_2 : _GEN_1215; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1217 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_2 : _GEN_1216; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1218 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_2 : _GEN_1217; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1219 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_2 : _GEN_1218; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1220 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_2 : _GEN_1219; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1221 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_2 : _GEN_1220; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1222 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_2 : _GEN_1221; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1223 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_2 : _GEN_1222; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1224 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_2 : _GEN_1223; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1225 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_2 : _GEN_1224; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1226 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_2 : _GEN_1225; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1227 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_2 : _GEN_1226; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1228 = dataModule_io_dataOut_0_2_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1229 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_5 : _GEN_1228; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1230 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_5 : _GEN_1229; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1231 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_5 : _GEN_1230; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1232 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_5 : _GEN_1231; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1233 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_5 : _GEN_1232; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1234 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_5 : _GEN_1233; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1235 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_5 : _GEN_1234; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1236 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_5 : _GEN_1235; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1237 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_5 : _GEN_1236; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1238 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_5 : _GEN_1237; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1239 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_5 : _GEN_1238; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1240 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_5 : _GEN_1239; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1241 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_5 : _GEN_1240; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1242 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_5 : _GEN_1241; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1243 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_5 : _GEN_1242; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1244 = dataModule_io_dataOut_0_2_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1245 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_4 : _GEN_1244; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1246 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_4 : _GEN_1245; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1247 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_4 : _GEN_1246; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1248 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_4 : _GEN_1247; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1249 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_4 : _GEN_1248; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1250 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_4 : _GEN_1249; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1251 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_4 : _GEN_1250; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1252 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_4 : _GEN_1251; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1253 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_4 : _GEN_1252; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1254 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_4 : _GEN_1253; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1255 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_4 : _GEN_1254; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1256 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_4 : _GEN_1255; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1257 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_4 : _GEN_1256; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1258 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_4 : _GEN_1257; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1259 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_4 : _GEN_1258; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1260 = dataModule_io_dataOut_0_2_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1261 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_7 : _GEN_1260; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1262 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_7 : _GEN_1261; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1263 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_7 : _GEN_1262; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1264 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_7 : _GEN_1263; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1265 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_7 : _GEN_1264; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1266 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_7 : _GEN_1265; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1267 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_7 : _GEN_1266; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1268 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_7 : _GEN_1267; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1269 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_7 : _GEN_1268; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1270 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_7 : _GEN_1269; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1271 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_7 : _GEN_1270; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1272 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_7 : _GEN_1271; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1273 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_7 : _GEN_1272; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1274 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_7 : _GEN_1273; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1275 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_7 : _GEN_1274; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1276 = dataModule_io_dataOut_0_2_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1277 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_2_6 : _GEN_1276; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1278 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_2_6 : _GEN_1277; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1279 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_2_6 : _GEN_1278; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1280 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_2_6 : _GEN_1279; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1281 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_2_6 : _GEN_1280; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1282 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_2_6 : _GEN_1281; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1283 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_2_6 : _GEN_1282; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1284 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_2_6 : _GEN_1283; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1285 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_2_6 : _GEN_1284; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1286 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_2_6 : _GEN_1285; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1287 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_2_6 : _GEN_1286; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1288 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_2_6 : _GEN_1287; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1289 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_2_6 : _GEN_1288; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1290 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_2_6 : _GEN_1289; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1291 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_2_6 : _GEN_1290; // @[Sbuffer.scala 703:{64,64}]
  wire [63:0] io_dcache_req_bits_data_lo_hi_lo = {_GEN_1275,_GEN_1291,_GEN_1243,_GEN_1259,_GEN_1211,_GEN_1227,_GEN_1179,
    _GEN_1195}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1292 = dataModule_io_dataOut_0_3_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1293 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_1 : _GEN_1292; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1294 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_1 : _GEN_1293; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1295 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_1 : _GEN_1294; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1296 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_1 : _GEN_1295; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1297 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_1 : _GEN_1296; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1298 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_1 : _GEN_1297; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1299 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_1 : _GEN_1298; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1300 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_1 : _GEN_1299; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1301 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_1 : _GEN_1300; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1302 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_1 : _GEN_1301; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1303 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_1 : _GEN_1302; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1304 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_1 : _GEN_1303; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1305 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_1 : _GEN_1304; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1306 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_1 : _GEN_1305; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1307 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_1 : _GEN_1306; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1308 = dataModule_io_dataOut_0_3_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1309 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_0 : _GEN_1308; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1310 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_0 : _GEN_1309; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1311 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_0 : _GEN_1310; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1312 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_0 : _GEN_1311; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1313 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_0 : _GEN_1312; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1314 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_0 : _GEN_1313; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1315 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_0 : _GEN_1314; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1316 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_0 : _GEN_1315; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1317 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_0 : _GEN_1316; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1318 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_0 : _GEN_1317; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1319 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_0 : _GEN_1318; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1320 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_0 : _GEN_1319; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1321 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_0 : _GEN_1320; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1322 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_0 : _GEN_1321; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1323 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_0 : _GEN_1322; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1324 = dataModule_io_dataOut_0_3_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1325 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_3 : _GEN_1324; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1326 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_3 : _GEN_1325; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1327 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_3 : _GEN_1326; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1328 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_3 : _GEN_1327; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1329 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_3 : _GEN_1328; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1330 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_3 : _GEN_1329; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1331 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_3 : _GEN_1330; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1332 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_3 : _GEN_1331; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1333 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_3 : _GEN_1332; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1334 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_3 : _GEN_1333; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1335 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_3 : _GEN_1334; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1336 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_3 : _GEN_1335; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1337 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_3 : _GEN_1336; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1338 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_3 : _GEN_1337; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1339 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_3 : _GEN_1338; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1340 = dataModule_io_dataOut_0_3_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1341 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_2 : _GEN_1340; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1342 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_2 : _GEN_1341; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1343 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_2 : _GEN_1342; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1344 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_2 : _GEN_1343; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1345 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_2 : _GEN_1344; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1346 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_2 : _GEN_1345; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1347 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_2 : _GEN_1346; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1348 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_2 : _GEN_1347; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1349 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_2 : _GEN_1348; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1350 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_2 : _GEN_1349; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1351 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_2 : _GEN_1350; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1352 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_2 : _GEN_1351; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1353 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_2 : _GEN_1352; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1354 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_2 : _GEN_1353; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1355 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_2 : _GEN_1354; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1356 = dataModule_io_dataOut_0_3_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1357 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_5 : _GEN_1356; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1358 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_5 : _GEN_1357; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1359 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_5 : _GEN_1358; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1360 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_5 : _GEN_1359; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1361 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_5 : _GEN_1360; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1362 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_5 : _GEN_1361; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1363 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_5 : _GEN_1362; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1364 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_5 : _GEN_1363; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1365 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_5 : _GEN_1364; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1366 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_5 : _GEN_1365; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1367 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_5 : _GEN_1366; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1368 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_5 : _GEN_1367; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1369 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_5 : _GEN_1368; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1370 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_5 : _GEN_1369; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1371 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_5 : _GEN_1370; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1372 = dataModule_io_dataOut_0_3_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1373 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_4 : _GEN_1372; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1374 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_4 : _GEN_1373; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1375 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_4 : _GEN_1374; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1376 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_4 : _GEN_1375; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1377 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_4 : _GEN_1376; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1378 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_4 : _GEN_1377; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1379 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_4 : _GEN_1378; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1380 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_4 : _GEN_1379; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1381 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_4 : _GEN_1380; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1382 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_4 : _GEN_1381; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1383 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_4 : _GEN_1382; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1384 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_4 : _GEN_1383; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1385 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_4 : _GEN_1384; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1386 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_4 : _GEN_1385; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1387 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_4 : _GEN_1386; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1388 = dataModule_io_dataOut_0_3_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1389 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_7 : _GEN_1388; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1390 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_7 : _GEN_1389; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1391 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_7 : _GEN_1390; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1392 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_7 : _GEN_1391; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1393 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_7 : _GEN_1392; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1394 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_7 : _GEN_1393; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1395 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_7 : _GEN_1394; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1396 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_7 : _GEN_1395; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1397 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_7 : _GEN_1396; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1398 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_7 : _GEN_1397; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1399 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_7 : _GEN_1398; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1400 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_7 : _GEN_1399; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1401 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_7 : _GEN_1400; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1402 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_7 : _GEN_1401; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1403 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_7 : _GEN_1402; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1404 = dataModule_io_dataOut_0_3_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1405 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_3_6 : _GEN_1404; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1406 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_3_6 : _GEN_1405; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1407 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_3_6 : _GEN_1406; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1408 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_3_6 : _GEN_1407; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1409 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_3_6 : _GEN_1408; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1410 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_3_6 : _GEN_1409; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1411 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_3_6 : _GEN_1410; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1412 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_3_6 : _GEN_1411; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1413 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_3_6 : _GEN_1412; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1414 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_3_6 : _GEN_1413; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1415 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_3_6 : _GEN_1414; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1416 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_3_6 : _GEN_1415; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1417 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_3_6 : _GEN_1416; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1418 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_3_6 : _GEN_1417; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1419 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_3_6 : _GEN_1418; // @[Sbuffer.scala 703:{64,64}]
  wire [255:0] io_dcache_req_bits_data_lo = {_GEN_1403,_GEN_1419,_GEN_1371,_GEN_1387,_GEN_1339,_GEN_1355,_GEN_1307,
    _GEN_1323,io_dcache_req_bits_data_lo_hi_lo,io_dcache_req_bits_data_lo_lo}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1420 = dataModule_io_dataOut_0_4_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1421 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_1 : _GEN_1420; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1422 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_1 : _GEN_1421; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1423 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_1 : _GEN_1422; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1424 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_1 : _GEN_1423; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1425 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_1 : _GEN_1424; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1426 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_1 : _GEN_1425; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1427 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_1 : _GEN_1426; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1428 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_1 : _GEN_1427; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1429 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_1 : _GEN_1428; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1430 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_1 : _GEN_1429; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1431 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_1 : _GEN_1430; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1432 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_1 : _GEN_1431; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1433 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_1 : _GEN_1432; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1434 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_1 : _GEN_1433; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1435 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_1 : _GEN_1434; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1436 = dataModule_io_dataOut_0_4_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1437 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_0 : _GEN_1436; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1438 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_0 : _GEN_1437; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1439 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_0 : _GEN_1438; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1440 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_0 : _GEN_1439; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1441 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_0 : _GEN_1440; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1442 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_0 : _GEN_1441; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1443 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_0 : _GEN_1442; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1444 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_0 : _GEN_1443; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1445 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_0 : _GEN_1444; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1446 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_0 : _GEN_1445; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1447 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_0 : _GEN_1446; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1448 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_0 : _GEN_1447; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1449 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_0 : _GEN_1448; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1450 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_0 : _GEN_1449; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1451 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_0 : _GEN_1450; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1452 = dataModule_io_dataOut_0_4_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1453 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_3 : _GEN_1452; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1454 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_3 : _GEN_1453; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1455 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_3 : _GEN_1454; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1456 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_3 : _GEN_1455; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1457 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_3 : _GEN_1456; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1458 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_3 : _GEN_1457; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1459 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_3 : _GEN_1458; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1460 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_3 : _GEN_1459; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1461 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_3 : _GEN_1460; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1462 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_3 : _GEN_1461; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1463 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_3 : _GEN_1462; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1464 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_3 : _GEN_1463; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1465 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_3 : _GEN_1464; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1466 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_3 : _GEN_1465; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1467 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_3 : _GEN_1466; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1468 = dataModule_io_dataOut_0_4_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1469 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_2 : _GEN_1468; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1470 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_2 : _GEN_1469; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1471 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_2 : _GEN_1470; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1472 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_2 : _GEN_1471; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1473 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_2 : _GEN_1472; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1474 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_2 : _GEN_1473; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1475 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_2 : _GEN_1474; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1476 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_2 : _GEN_1475; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1477 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_2 : _GEN_1476; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1478 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_2 : _GEN_1477; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1479 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_2 : _GEN_1478; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1480 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_2 : _GEN_1479; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1481 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_2 : _GEN_1480; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1482 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_2 : _GEN_1481; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1483 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_2 : _GEN_1482; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1484 = dataModule_io_dataOut_0_4_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1485 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_5 : _GEN_1484; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1486 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_5 : _GEN_1485; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1487 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_5 : _GEN_1486; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1488 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_5 : _GEN_1487; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1489 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_5 : _GEN_1488; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1490 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_5 : _GEN_1489; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1491 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_5 : _GEN_1490; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1492 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_5 : _GEN_1491; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1493 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_5 : _GEN_1492; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1494 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_5 : _GEN_1493; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1495 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_5 : _GEN_1494; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1496 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_5 : _GEN_1495; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1497 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_5 : _GEN_1496; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1498 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_5 : _GEN_1497; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1499 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_5 : _GEN_1498; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1500 = dataModule_io_dataOut_0_4_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1501 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_4 : _GEN_1500; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1502 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_4 : _GEN_1501; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1503 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_4 : _GEN_1502; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1504 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_4 : _GEN_1503; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1505 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_4 : _GEN_1504; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1506 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_4 : _GEN_1505; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1507 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_4 : _GEN_1506; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1508 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_4 : _GEN_1507; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1509 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_4 : _GEN_1508; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1510 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_4 : _GEN_1509; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1511 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_4 : _GEN_1510; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1512 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_4 : _GEN_1511; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1513 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_4 : _GEN_1512; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1514 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_4 : _GEN_1513; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1515 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_4 : _GEN_1514; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1516 = dataModule_io_dataOut_0_4_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1517 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_7 : _GEN_1516; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1518 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_7 : _GEN_1517; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1519 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_7 : _GEN_1518; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1520 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_7 : _GEN_1519; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1521 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_7 : _GEN_1520; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1522 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_7 : _GEN_1521; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1523 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_7 : _GEN_1522; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1524 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_7 : _GEN_1523; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1525 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_7 : _GEN_1524; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1526 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_7 : _GEN_1525; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1527 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_7 : _GEN_1526; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1528 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_7 : _GEN_1527; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1529 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_7 : _GEN_1528; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1530 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_7 : _GEN_1529; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1531 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_7 : _GEN_1530; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1532 = dataModule_io_dataOut_0_4_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1533 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_4_6 : _GEN_1532; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1534 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_4_6 : _GEN_1533; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1535 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_4_6 : _GEN_1534; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1536 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_4_6 : _GEN_1535; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1537 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_4_6 : _GEN_1536; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1538 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_4_6 : _GEN_1537; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1539 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_4_6 : _GEN_1538; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1540 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_4_6 : _GEN_1539; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1541 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_4_6 : _GEN_1540; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1542 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_4_6 : _GEN_1541; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1543 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_4_6 : _GEN_1542; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1544 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_4_6 : _GEN_1543; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1545 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_4_6 : _GEN_1544; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1546 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_4_6 : _GEN_1545; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1547 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_4_6 : _GEN_1546; // @[Sbuffer.scala 703:{64,64}]
  wire [63:0] io_dcache_req_bits_data_hi_lo_lo = {_GEN_1531,_GEN_1547,_GEN_1499,_GEN_1515,_GEN_1467,_GEN_1483,_GEN_1435,
    _GEN_1451}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1548 = dataModule_io_dataOut_0_5_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1549 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_1 : _GEN_1548; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1550 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_1 : _GEN_1549; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1551 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_1 : _GEN_1550; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1552 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_1 : _GEN_1551; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1553 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_1 : _GEN_1552; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1554 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_1 : _GEN_1553; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1555 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_1 : _GEN_1554; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1556 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_1 : _GEN_1555; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1557 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_1 : _GEN_1556; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1558 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_1 : _GEN_1557; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1559 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_1 : _GEN_1558; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1560 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_1 : _GEN_1559; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1561 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_1 : _GEN_1560; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1562 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_1 : _GEN_1561; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1563 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_1 : _GEN_1562; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1564 = dataModule_io_dataOut_0_5_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1565 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_0 : _GEN_1564; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1566 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_0 : _GEN_1565; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1567 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_0 : _GEN_1566; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1568 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_0 : _GEN_1567; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1569 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_0 : _GEN_1568; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1570 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_0 : _GEN_1569; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1571 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_0 : _GEN_1570; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1572 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_0 : _GEN_1571; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1573 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_0 : _GEN_1572; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1574 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_0 : _GEN_1573; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1575 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_0 : _GEN_1574; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1576 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_0 : _GEN_1575; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1577 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_0 : _GEN_1576; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1578 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_0 : _GEN_1577; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1579 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_0 : _GEN_1578; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1580 = dataModule_io_dataOut_0_5_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1581 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_3 : _GEN_1580; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1582 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_3 : _GEN_1581; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1583 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_3 : _GEN_1582; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1584 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_3 : _GEN_1583; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1585 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_3 : _GEN_1584; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1586 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_3 : _GEN_1585; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1587 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_3 : _GEN_1586; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1588 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_3 : _GEN_1587; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1589 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_3 : _GEN_1588; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1590 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_3 : _GEN_1589; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1591 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_3 : _GEN_1590; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1592 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_3 : _GEN_1591; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1593 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_3 : _GEN_1592; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1594 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_3 : _GEN_1593; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1595 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_3 : _GEN_1594; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1596 = dataModule_io_dataOut_0_5_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1597 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_2 : _GEN_1596; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1598 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_2 : _GEN_1597; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1599 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_2 : _GEN_1598; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1600 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_2 : _GEN_1599; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1601 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_2 : _GEN_1600; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1602 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_2 : _GEN_1601; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1603 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_2 : _GEN_1602; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1604 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_2 : _GEN_1603; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1605 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_2 : _GEN_1604; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1606 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_2 : _GEN_1605; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1607 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_2 : _GEN_1606; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1608 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_2 : _GEN_1607; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1609 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_2 : _GEN_1608; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1610 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_2 : _GEN_1609; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1611 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_2 : _GEN_1610; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1612 = dataModule_io_dataOut_0_5_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1613 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_5 : _GEN_1612; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1614 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_5 : _GEN_1613; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1615 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_5 : _GEN_1614; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1616 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_5 : _GEN_1615; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1617 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_5 : _GEN_1616; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1618 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_5 : _GEN_1617; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1619 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_5 : _GEN_1618; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1620 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_5 : _GEN_1619; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1621 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_5 : _GEN_1620; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1622 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_5 : _GEN_1621; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1623 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_5 : _GEN_1622; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1624 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_5 : _GEN_1623; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1625 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_5 : _GEN_1624; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1626 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_5 : _GEN_1625; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1627 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_5 : _GEN_1626; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1628 = dataModule_io_dataOut_0_5_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1629 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_4 : _GEN_1628; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1630 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_4 : _GEN_1629; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1631 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_4 : _GEN_1630; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1632 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_4 : _GEN_1631; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1633 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_4 : _GEN_1632; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1634 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_4 : _GEN_1633; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1635 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_4 : _GEN_1634; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1636 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_4 : _GEN_1635; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1637 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_4 : _GEN_1636; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1638 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_4 : _GEN_1637; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1639 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_4 : _GEN_1638; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1640 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_4 : _GEN_1639; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1641 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_4 : _GEN_1640; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1642 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_4 : _GEN_1641; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1643 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_4 : _GEN_1642; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1644 = dataModule_io_dataOut_0_5_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1645 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_7 : _GEN_1644; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1646 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_7 : _GEN_1645; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1647 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_7 : _GEN_1646; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1648 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_7 : _GEN_1647; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1649 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_7 : _GEN_1648; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1650 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_7 : _GEN_1649; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1651 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_7 : _GEN_1650; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1652 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_7 : _GEN_1651; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1653 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_7 : _GEN_1652; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1654 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_7 : _GEN_1653; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1655 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_7 : _GEN_1654; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1656 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_7 : _GEN_1655; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1657 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_7 : _GEN_1656; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1658 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_7 : _GEN_1657; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1659 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_7 : _GEN_1658; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1660 = dataModule_io_dataOut_0_5_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1661 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_5_6 : _GEN_1660; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1662 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_5_6 : _GEN_1661; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1663 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_5_6 : _GEN_1662; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1664 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_5_6 : _GEN_1663; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1665 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_5_6 : _GEN_1664; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1666 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_5_6 : _GEN_1665; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1667 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_5_6 : _GEN_1666; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1668 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_5_6 : _GEN_1667; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1669 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_5_6 : _GEN_1668; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1670 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_5_6 : _GEN_1669; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1671 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_5_6 : _GEN_1670; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1672 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_5_6 : _GEN_1671; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1673 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_5_6 : _GEN_1672; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1674 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_5_6 : _GEN_1673; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1675 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_5_6 : _GEN_1674; // @[Sbuffer.scala 703:{64,64}]
  wire [127:0] io_dcache_req_bits_data_hi_lo = {_GEN_1659,_GEN_1675,_GEN_1627,_GEN_1643,_GEN_1595,_GEN_1611,_GEN_1563,
    _GEN_1579,io_dcache_req_bits_data_hi_lo_lo}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1676 = dataModule_io_dataOut_0_6_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1677 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_1 : _GEN_1676; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1678 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_1 : _GEN_1677; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1679 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_1 : _GEN_1678; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1680 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_1 : _GEN_1679; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1681 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_1 : _GEN_1680; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1682 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_1 : _GEN_1681; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1683 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_1 : _GEN_1682; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1684 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_1 : _GEN_1683; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1685 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_1 : _GEN_1684; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1686 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_1 : _GEN_1685; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1687 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_1 : _GEN_1686; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1688 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_1 : _GEN_1687; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1689 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_1 : _GEN_1688; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1690 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_1 : _GEN_1689; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1691 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_1 : _GEN_1690; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1692 = dataModule_io_dataOut_0_6_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1693 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_0 : _GEN_1692; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1694 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_0 : _GEN_1693; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1695 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_0 : _GEN_1694; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1696 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_0 : _GEN_1695; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1697 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_0 : _GEN_1696; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1698 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_0 : _GEN_1697; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1699 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_0 : _GEN_1698; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1700 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_0 : _GEN_1699; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1701 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_0 : _GEN_1700; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1702 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_0 : _GEN_1701; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1703 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_0 : _GEN_1702; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1704 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_0 : _GEN_1703; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1705 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_0 : _GEN_1704; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1706 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_0 : _GEN_1705; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1707 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_0 : _GEN_1706; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1708 = dataModule_io_dataOut_0_6_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1709 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_3 : _GEN_1708; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1710 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_3 : _GEN_1709; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1711 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_3 : _GEN_1710; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1712 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_3 : _GEN_1711; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1713 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_3 : _GEN_1712; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1714 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_3 : _GEN_1713; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1715 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_3 : _GEN_1714; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1716 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_3 : _GEN_1715; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1717 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_3 : _GEN_1716; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1718 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_3 : _GEN_1717; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1719 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_3 : _GEN_1718; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1720 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_3 : _GEN_1719; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1721 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_3 : _GEN_1720; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1722 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_3 : _GEN_1721; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1723 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_3 : _GEN_1722; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1724 = dataModule_io_dataOut_0_6_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1725 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_2 : _GEN_1724; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1726 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_2 : _GEN_1725; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1727 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_2 : _GEN_1726; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1728 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_2 : _GEN_1727; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1729 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_2 : _GEN_1728; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1730 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_2 : _GEN_1729; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1731 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_2 : _GEN_1730; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1732 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_2 : _GEN_1731; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1733 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_2 : _GEN_1732; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1734 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_2 : _GEN_1733; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1735 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_2 : _GEN_1734; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1736 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_2 : _GEN_1735; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1737 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_2 : _GEN_1736; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1738 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_2 : _GEN_1737; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1739 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_2 : _GEN_1738; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1740 = dataModule_io_dataOut_0_6_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1741 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_5 : _GEN_1740; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1742 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_5 : _GEN_1741; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1743 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_5 : _GEN_1742; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1744 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_5 : _GEN_1743; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1745 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_5 : _GEN_1744; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1746 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_5 : _GEN_1745; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1747 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_5 : _GEN_1746; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1748 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_5 : _GEN_1747; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1749 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_5 : _GEN_1748; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1750 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_5 : _GEN_1749; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1751 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_5 : _GEN_1750; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1752 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_5 : _GEN_1751; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1753 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_5 : _GEN_1752; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1754 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_5 : _GEN_1753; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1755 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_5 : _GEN_1754; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1756 = dataModule_io_dataOut_0_6_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1757 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_4 : _GEN_1756; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1758 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_4 : _GEN_1757; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1759 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_4 : _GEN_1758; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1760 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_4 : _GEN_1759; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1761 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_4 : _GEN_1760; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1762 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_4 : _GEN_1761; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1763 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_4 : _GEN_1762; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1764 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_4 : _GEN_1763; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1765 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_4 : _GEN_1764; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1766 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_4 : _GEN_1765; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1767 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_4 : _GEN_1766; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1768 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_4 : _GEN_1767; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1769 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_4 : _GEN_1768; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1770 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_4 : _GEN_1769; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1771 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_4 : _GEN_1770; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1772 = dataModule_io_dataOut_0_6_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1773 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_7 : _GEN_1772; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1774 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_7 : _GEN_1773; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1775 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_7 : _GEN_1774; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1776 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_7 : _GEN_1775; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1777 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_7 : _GEN_1776; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1778 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_7 : _GEN_1777; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1779 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_7 : _GEN_1778; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1780 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_7 : _GEN_1779; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1781 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_7 : _GEN_1780; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1782 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_7 : _GEN_1781; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1783 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_7 : _GEN_1782; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1784 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_7 : _GEN_1783; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1785 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_7 : _GEN_1784; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1786 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_7 : _GEN_1785; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1787 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_7 : _GEN_1786; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1788 = dataModule_io_dataOut_0_6_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1789 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_6_6 : _GEN_1788; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1790 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_6_6 : _GEN_1789; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1791 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_6_6 : _GEN_1790; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1792 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_6_6 : _GEN_1791; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1793 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_6_6 : _GEN_1792; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1794 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_6_6 : _GEN_1793; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1795 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_6_6 : _GEN_1794; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1796 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_6_6 : _GEN_1795; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1797 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_6_6 : _GEN_1796; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1798 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_6_6 : _GEN_1797; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1799 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_6_6 : _GEN_1798; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1800 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_6_6 : _GEN_1799; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1801 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_6_6 : _GEN_1800; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1802 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_6_6 : _GEN_1801; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1803 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_6_6 : _GEN_1802; // @[Sbuffer.scala 703:{64,64}]
  wire [63:0] io_dcache_req_bits_data_hi_hi_lo = {_GEN_1787,_GEN_1803,_GEN_1755,_GEN_1771,_GEN_1723,_GEN_1739,_GEN_1691,
    _GEN_1707}; // @[Sbuffer.scala 703:64]
  wire [7:0] _GEN_1804 = dataModule_io_dataOut_0_7_1; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1805 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_1 : _GEN_1804; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1806 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_1 : _GEN_1805; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1807 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_1 : _GEN_1806; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1808 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_1 : _GEN_1807; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1809 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_1 : _GEN_1808; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1810 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_1 : _GEN_1809; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1811 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_1 : _GEN_1810; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1812 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_1 : _GEN_1811; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1813 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_1 : _GEN_1812; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1814 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_1 : _GEN_1813; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1815 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_1 : _GEN_1814; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1816 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_1 : _GEN_1815; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1817 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_1 : _GEN_1816; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1818 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_1 : _GEN_1817; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1819 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_1 : _GEN_1818; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1820 = dataModule_io_dataOut_0_7_0; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1821 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_0 : _GEN_1820; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1822 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_0 : _GEN_1821; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1823 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_0 : _GEN_1822; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1824 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_0 : _GEN_1823; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1825 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_0 : _GEN_1824; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1826 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_0 : _GEN_1825; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1827 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_0 : _GEN_1826; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1828 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_0 : _GEN_1827; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1829 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_0 : _GEN_1828; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1830 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_0 : _GEN_1829; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1831 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_0 : _GEN_1830; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1832 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_0 : _GEN_1831; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1833 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_0 : _GEN_1832; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1834 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_0 : _GEN_1833; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1835 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_0 : _GEN_1834; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1836 = dataModule_io_dataOut_0_7_3; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1837 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_3 : _GEN_1836; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1838 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_3 : _GEN_1837; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1839 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_3 : _GEN_1838; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1840 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_3 : _GEN_1839; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1841 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_3 : _GEN_1840; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1842 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_3 : _GEN_1841; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1843 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_3 : _GEN_1842; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1844 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_3 : _GEN_1843; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1845 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_3 : _GEN_1844; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1846 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_3 : _GEN_1845; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1847 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_3 : _GEN_1846; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1848 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_3 : _GEN_1847; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1849 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_3 : _GEN_1848; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1850 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_3 : _GEN_1849; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1851 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_3 : _GEN_1850; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1852 = dataModule_io_dataOut_0_7_2; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1853 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_2 : _GEN_1852; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1854 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_2 : _GEN_1853; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1855 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_2 : _GEN_1854; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1856 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_2 : _GEN_1855; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1857 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_2 : _GEN_1856; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1858 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_2 : _GEN_1857; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1859 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_2 : _GEN_1858; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1860 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_2 : _GEN_1859; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1861 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_2 : _GEN_1860; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1862 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_2 : _GEN_1861; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1863 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_2 : _GEN_1862; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1864 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_2 : _GEN_1863; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1865 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_2 : _GEN_1864; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1866 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_2 : _GEN_1865; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1867 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_2 : _GEN_1866; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1868 = dataModule_io_dataOut_0_7_5; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1869 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_5 : _GEN_1868; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1870 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_5 : _GEN_1869; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1871 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_5 : _GEN_1870; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1872 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_5 : _GEN_1871; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1873 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_5 : _GEN_1872; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1874 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_5 : _GEN_1873; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1875 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_5 : _GEN_1874; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1876 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_5 : _GEN_1875; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1877 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_5 : _GEN_1876; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1878 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_5 : _GEN_1877; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1879 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_5 : _GEN_1878; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1880 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_5 : _GEN_1879; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1881 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_5 : _GEN_1880; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1882 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_5 : _GEN_1881; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1883 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_5 : _GEN_1882; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1884 = dataModule_io_dataOut_0_7_4; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1885 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_4 : _GEN_1884; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1886 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_4 : _GEN_1885; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1887 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_4 : _GEN_1886; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1888 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_4 : _GEN_1887; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1889 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_4 : _GEN_1888; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1890 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_4 : _GEN_1889; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1891 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_4 : _GEN_1890; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1892 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_4 : _GEN_1891; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1893 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_4 : _GEN_1892; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1894 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_4 : _GEN_1893; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1895 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_4 : _GEN_1894; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1896 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_4 : _GEN_1895; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1897 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_4 : _GEN_1896; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1898 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_4 : _GEN_1897; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1899 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_4 : _GEN_1898; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1900 = dataModule_io_dataOut_0_7_7; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1901 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_7 : _GEN_1900; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1902 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_7 : _GEN_1901; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1903 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_7 : _GEN_1902; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1904 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_7 : _GEN_1903; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1905 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_7 : _GEN_1904; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1906 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_7 : _GEN_1905; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1907 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_7 : _GEN_1906; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1908 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_7 : _GEN_1907; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1909 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_7 : _GEN_1908; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1910 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_7 : _GEN_1909; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1911 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_7 : _GEN_1910; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1912 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_7 : _GEN_1911; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1913 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_7 : _GEN_1912; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1914 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_7 : _GEN_1913; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1915 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_7 : _GEN_1914; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1916 = dataModule_io_dataOut_0_7_6; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1917 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_1_7_6 : _GEN_1916; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1918 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_2_7_6 : _GEN_1917; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1919 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_3_7_6 : _GEN_1918; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1920 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_4_7_6 : _GEN_1919; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1921 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_5_7_6 : _GEN_1920; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1922 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_6_7_6 : _GEN_1921; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1923 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_7_7_6 : _GEN_1922; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1924 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_8_7_6 : _GEN_1923; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1925 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_9_7_6 : _GEN_1924; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1926 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_10_7_6 : _GEN_1925; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1927 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_11_7_6 : _GEN_1926; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1928 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_12_7_6 : _GEN_1927; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1929 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_13_7_6 : _GEN_1928; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1930 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_14_7_6 : _GEN_1929; // @[Sbuffer.scala 703:{64,64}]
  wire [7:0] _GEN_1931 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_dataOut_15_7_6 : _GEN_1930; // @[Sbuffer.scala 703:{64,64}]
  wire [255:0] io_dcache_req_bits_data_hi = {_GEN_1915,_GEN_1931,_GEN_1883,_GEN_1899,_GEN_1851,_GEN_1867,_GEN_1819,
    _GEN_1835,io_dcache_req_bits_data_hi_hi_lo,io_dcache_req_bits_data_hi_lo}; // @[Sbuffer.scala 703:64]
  wire  _GEN_1932 = dataModule_io_maskOut_0_0_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1933 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_1 : dataModule_io_maskOut_0_0_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1934 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_1 : _GEN_1933; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1935 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_1 : _GEN_1934; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1936 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_1 : _GEN_1935; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1937 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_1 : _GEN_1936; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1938 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_1 : _GEN_1937; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1939 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_1 : _GEN_1938; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1940 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_1 : _GEN_1939; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1941 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_1 : _GEN_1940; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1942 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_1 : _GEN_1941; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1943 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_1 : _GEN_1942; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1944 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_1 : _GEN_1943; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1945 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_1 : _GEN_1944; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1946 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_1 : _GEN_1945; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1947 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_1 : _GEN_1946; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1948 = dataModule_io_maskOut_0_0_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1949 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_0 : dataModule_io_maskOut_0_0_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1950 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_0 : _GEN_1949; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1951 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_0 : _GEN_1950; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1952 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_0 : _GEN_1951; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1953 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_0 : _GEN_1952; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1954 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_0 : _GEN_1953; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1955 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_0 : _GEN_1954; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1956 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_0 : _GEN_1955; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1957 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_0 : _GEN_1956; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1958 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_0 : _GEN_1957; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1959 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_0 : _GEN_1958; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1960 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_0 : _GEN_1959; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1961 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_0 : _GEN_1960; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1962 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_0 : _GEN_1961; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1963 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_0 : _GEN_1962; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1964 = dataModule_io_maskOut_0_0_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1965 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_3 : dataModule_io_maskOut_0_0_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1966 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_3 : _GEN_1965; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1967 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_3 : _GEN_1966; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1968 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_3 : _GEN_1967; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1969 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_3 : _GEN_1968; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1970 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_3 : _GEN_1969; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1971 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_3 : _GEN_1970; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1972 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_3 : _GEN_1971; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1973 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_3 : _GEN_1972; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1974 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_3 : _GEN_1973; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1975 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_3 : _GEN_1974; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1976 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_3 : _GEN_1975; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1977 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_3 : _GEN_1976; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1978 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_3 : _GEN_1977; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1979 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_3 : _GEN_1978; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1980 = dataModule_io_maskOut_0_0_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1981 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_2 : dataModule_io_maskOut_0_0_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1982 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_2 : _GEN_1981; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1983 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_2 : _GEN_1982; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1984 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_2 : _GEN_1983; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1985 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_2 : _GEN_1984; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1986 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_2 : _GEN_1985; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1987 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_2 : _GEN_1986; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1988 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_2 : _GEN_1987; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1989 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_2 : _GEN_1988; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1990 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_2 : _GEN_1989; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1991 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_2 : _GEN_1990; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1992 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_2 : _GEN_1991; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1993 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_2 : _GEN_1992; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1994 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_2 : _GEN_1993; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1995 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_2 : _GEN_1994; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1996 = dataModule_io_maskOut_0_0_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1997 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_5 : dataModule_io_maskOut_0_0_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1998 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_5 : _GEN_1997; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_1999 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_5 : _GEN_1998; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2000 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_5 : _GEN_1999; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2001 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_5 : _GEN_2000; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2002 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_5 : _GEN_2001; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2003 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_5 : _GEN_2002; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2004 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_5 : _GEN_2003; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2005 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_5 : _GEN_2004; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2006 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_5 : _GEN_2005; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2007 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_5 : _GEN_2006; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2008 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_5 : _GEN_2007; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2009 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_5 : _GEN_2008; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2010 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_5 : _GEN_2009; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2011 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_5 : _GEN_2010; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2012 = dataModule_io_maskOut_0_0_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2013 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_4 : dataModule_io_maskOut_0_0_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2014 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_4 : _GEN_2013; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2015 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_4 : _GEN_2014; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2016 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_4 : _GEN_2015; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2017 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_4 : _GEN_2016; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2018 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_4 : _GEN_2017; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2019 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_4 : _GEN_2018; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2020 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_4 : _GEN_2019; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2021 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_4 : _GEN_2020; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2022 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_4 : _GEN_2021; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2023 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_4 : _GEN_2022; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2024 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_4 : _GEN_2023; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2025 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_4 : _GEN_2024; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2026 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_4 : _GEN_2025; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2027 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_4 : _GEN_2026; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2028 = dataModule_io_maskOut_0_0_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2029 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_7 : dataModule_io_maskOut_0_0_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2030 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_7 : _GEN_2029; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2031 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_7 : _GEN_2030; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2032 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_7 : _GEN_2031; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2033 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_7 : _GEN_2032; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2034 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_7 : _GEN_2033; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2035 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_7 : _GEN_2034; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2036 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_7 : _GEN_2035; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2037 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_7 : _GEN_2036; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2038 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_7 : _GEN_2037; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2039 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_7 : _GEN_2038; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2040 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_7 : _GEN_2039; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2041 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_7 : _GEN_2040; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2042 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_7 : _GEN_2041; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2043 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_7 : _GEN_2042; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2044 = dataModule_io_maskOut_0_0_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2045 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_0_6 : dataModule_io_maskOut_0_0_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2046 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_0_6 : _GEN_2045; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2047 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_0_6 : _GEN_2046; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2048 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_0_6 : _GEN_2047; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2049 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_0_6 : _GEN_2048; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2050 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_0_6 : _GEN_2049; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2051 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_0_6 : _GEN_2050; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2052 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_0_6 : _GEN_2051; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2053 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_0_6 : _GEN_2052; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2054 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_0_6 : _GEN_2053; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2055 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_0_6 : _GEN_2054; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2056 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_0_6 : _GEN_2055; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2057 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_0_6 : _GEN_2056; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2058 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_0_6 : _GEN_2057; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2059 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_0_6 : _GEN_2058; // @[Sbuffer.scala 704:{64,64}]
  wire [7:0] io_dcache_req_bits_mask_lo_lo_lo = {_GEN_2043,_GEN_2059,_GEN_2011,_GEN_2027,_GEN_1979,_GEN_1995,_GEN_1947,
    _GEN_1963}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2061 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_1 : dataModule_io_maskOut_0_1_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2062 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_1 : _GEN_2061; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2063 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_1 : _GEN_2062; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2064 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_1 : _GEN_2063; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2065 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_1 : _GEN_2064; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2066 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_1 : _GEN_2065; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2067 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_1 : _GEN_2066; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2068 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_1 : _GEN_2067; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2069 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_1 : _GEN_2068; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2070 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_1 : _GEN_2069; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2071 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_1 : _GEN_2070; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2072 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_1 : _GEN_2071; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2073 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_1 : _GEN_2072; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2074 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_1 : _GEN_2073; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2075 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_1 : _GEN_2074; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2077 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_0 : dataModule_io_maskOut_0_1_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2078 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_0 : _GEN_2077; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2079 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_0 : _GEN_2078; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2080 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_0 : _GEN_2079; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2081 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_0 : _GEN_2080; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2082 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_0 : _GEN_2081; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2083 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_0 : _GEN_2082; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2084 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_0 : _GEN_2083; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2085 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_0 : _GEN_2084; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2086 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_0 : _GEN_2085; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2087 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_0 : _GEN_2086; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2088 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_0 : _GEN_2087; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2089 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_0 : _GEN_2088; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2090 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_0 : _GEN_2089; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2091 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_0 : _GEN_2090; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2093 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_3 : dataModule_io_maskOut_0_1_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2094 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_3 : _GEN_2093; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2095 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_3 : _GEN_2094; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2096 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_3 : _GEN_2095; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2097 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_3 : _GEN_2096; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2098 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_3 : _GEN_2097; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2099 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_3 : _GEN_2098; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2100 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_3 : _GEN_2099; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2101 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_3 : _GEN_2100; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2102 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_3 : _GEN_2101; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2103 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_3 : _GEN_2102; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2104 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_3 : _GEN_2103; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2105 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_3 : _GEN_2104; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2106 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_3 : _GEN_2105; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2107 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_3 : _GEN_2106; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2109 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_2 : dataModule_io_maskOut_0_1_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2110 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_2 : _GEN_2109; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2111 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_2 : _GEN_2110; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2112 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_2 : _GEN_2111; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2113 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_2 : _GEN_2112; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2114 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_2 : _GEN_2113; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2115 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_2 : _GEN_2114; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2116 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_2 : _GEN_2115; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2117 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_2 : _GEN_2116; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2118 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_2 : _GEN_2117; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2119 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_2 : _GEN_2118; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2120 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_2 : _GEN_2119; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2121 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_2 : _GEN_2120; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2122 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_2 : _GEN_2121; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2123 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_2 : _GEN_2122; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2125 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_5 : dataModule_io_maskOut_0_1_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2126 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_5 : _GEN_2125; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2127 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_5 : _GEN_2126; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2128 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_5 : _GEN_2127; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2129 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_5 : _GEN_2128; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2130 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_5 : _GEN_2129; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2131 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_5 : _GEN_2130; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2132 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_5 : _GEN_2131; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2133 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_5 : _GEN_2132; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2134 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_5 : _GEN_2133; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2135 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_5 : _GEN_2134; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2136 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_5 : _GEN_2135; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2137 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_5 : _GEN_2136; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2138 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_5 : _GEN_2137; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2139 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_5 : _GEN_2138; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2141 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_4 : dataModule_io_maskOut_0_1_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2142 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_4 : _GEN_2141; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2143 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_4 : _GEN_2142; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2144 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_4 : _GEN_2143; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2145 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_4 : _GEN_2144; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2146 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_4 : _GEN_2145; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2147 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_4 : _GEN_2146; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2148 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_4 : _GEN_2147; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2149 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_4 : _GEN_2148; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2150 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_4 : _GEN_2149; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2151 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_4 : _GEN_2150; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2152 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_4 : _GEN_2151; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2153 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_4 : _GEN_2152; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2154 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_4 : _GEN_2153; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2155 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_4 : _GEN_2154; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2157 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_7 : dataModule_io_maskOut_0_1_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2158 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_7 : _GEN_2157; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2159 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_7 : _GEN_2158; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2160 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_7 : _GEN_2159; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2161 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_7 : _GEN_2160; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2162 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_7 : _GEN_2161; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2163 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_7 : _GEN_2162; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2164 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_7 : _GEN_2163; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2165 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_7 : _GEN_2164; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2166 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_7 : _GEN_2165; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2167 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_7 : _GEN_2166; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2168 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_7 : _GEN_2167; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2169 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_7 : _GEN_2168; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2170 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_7 : _GEN_2169; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2171 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_7 : _GEN_2170; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2173 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_1_6 : dataModule_io_maskOut_0_1_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2174 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_1_6 : _GEN_2173; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2175 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_1_6 : _GEN_2174; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2176 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_1_6 : _GEN_2175; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2177 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_1_6 : _GEN_2176; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2178 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_1_6 : _GEN_2177; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2179 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_1_6 : _GEN_2178; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2180 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_1_6 : _GEN_2179; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2181 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_1_6 : _GEN_2180; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2182 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_1_6 : _GEN_2181; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2183 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_1_6 : _GEN_2182; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2184 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_1_6 : _GEN_2183; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2185 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_1_6 : _GEN_2184; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2186 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_1_6 : _GEN_2185; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2187 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_1_6 : _GEN_2186; // @[Sbuffer.scala 704:{64,64}]
  wire [15:0] io_dcache_req_bits_mask_lo_lo = {_GEN_2171,_GEN_2187,_GEN_2139,_GEN_2155,_GEN_2107,_GEN_2123,_GEN_2075,
    _GEN_2091,io_dcache_req_bits_mask_lo_lo_lo}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2189 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_1 : dataModule_io_maskOut_0_2_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2190 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_1 : _GEN_2189; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2191 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_1 : _GEN_2190; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2192 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_1 : _GEN_2191; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2193 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_1 : _GEN_2192; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2194 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_1 : _GEN_2193; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2195 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_1 : _GEN_2194; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2196 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_1 : _GEN_2195; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2197 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_1 : _GEN_2196; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2198 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_1 : _GEN_2197; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2199 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_1 : _GEN_2198; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2200 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_1 : _GEN_2199; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2201 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_1 : _GEN_2200; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2202 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_1 : _GEN_2201; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2203 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_1 : _GEN_2202; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2205 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_0 : dataModule_io_maskOut_0_2_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2206 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_0 : _GEN_2205; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2207 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_0 : _GEN_2206; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2208 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_0 : _GEN_2207; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2209 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_0 : _GEN_2208; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2210 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_0 : _GEN_2209; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2211 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_0 : _GEN_2210; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2212 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_0 : _GEN_2211; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2213 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_0 : _GEN_2212; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2214 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_0 : _GEN_2213; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2215 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_0 : _GEN_2214; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2216 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_0 : _GEN_2215; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2217 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_0 : _GEN_2216; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2218 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_0 : _GEN_2217; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2219 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_0 : _GEN_2218; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2221 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_3 : dataModule_io_maskOut_0_2_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2222 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_3 : _GEN_2221; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2223 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_3 : _GEN_2222; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2224 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_3 : _GEN_2223; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2225 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_3 : _GEN_2224; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2226 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_3 : _GEN_2225; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2227 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_3 : _GEN_2226; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2228 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_3 : _GEN_2227; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2229 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_3 : _GEN_2228; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2230 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_3 : _GEN_2229; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2231 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_3 : _GEN_2230; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2232 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_3 : _GEN_2231; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2233 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_3 : _GEN_2232; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2234 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_3 : _GEN_2233; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2235 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_3 : _GEN_2234; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2237 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_2 : dataModule_io_maskOut_0_2_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2238 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_2 : _GEN_2237; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2239 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_2 : _GEN_2238; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2240 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_2 : _GEN_2239; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2241 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_2 : _GEN_2240; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2242 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_2 : _GEN_2241; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2243 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_2 : _GEN_2242; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2244 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_2 : _GEN_2243; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2245 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_2 : _GEN_2244; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2246 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_2 : _GEN_2245; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2247 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_2 : _GEN_2246; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2248 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_2 : _GEN_2247; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2249 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_2 : _GEN_2248; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2250 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_2 : _GEN_2249; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2251 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_2 : _GEN_2250; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2253 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_5 : dataModule_io_maskOut_0_2_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2254 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_5 : _GEN_2253; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2255 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_5 : _GEN_2254; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2256 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_5 : _GEN_2255; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2257 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_5 : _GEN_2256; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2258 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_5 : _GEN_2257; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2259 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_5 : _GEN_2258; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2260 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_5 : _GEN_2259; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2261 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_5 : _GEN_2260; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2262 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_5 : _GEN_2261; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2263 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_5 : _GEN_2262; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2264 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_5 : _GEN_2263; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2265 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_5 : _GEN_2264; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2266 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_5 : _GEN_2265; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2267 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_5 : _GEN_2266; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2269 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_4 : dataModule_io_maskOut_0_2_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2270 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_4 : _GEN_2269; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2271 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_4 : _GEN_2270; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2272 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_4 : _GEN_2271; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2273 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_4 : _GEN_2272; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2274 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_4 : _GEN_2273; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2275 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_4 : _GEN_2274; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2276 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_4 : _GEN_2275; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2277 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_4 : _GEN_2276; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2278 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_4 : _GEN_2277; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2279 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_4 : _GEN_2278; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2280 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_4 : _GEN_2279; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2281 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_4 : _GEN_2280; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2282 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_4 : _GEN_2281; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2283 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_4 : _GEN_2282; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2285 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_7 : dataModule_io_maskOut_0_2_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2286 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_7 : _GEN_2285; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2287 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_7 : _GEN_2286; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2288 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_7 : _GEN_2287; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2289 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_7 : _GEN_2288; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2290 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_7 : _GEN_2289; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2291 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_7 : _GEN_2290; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2292 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_7 : _GEN_2291; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2293 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_7 : _GEN_2292; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2294 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_7 : _GEN_2293; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2295 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_7 : _GEN_2294; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2296 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_7 : _GEN_2295; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2297 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_7 : _GEN_2296; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2298 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_7 : _GEN_2297; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2299 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_7 : _GEN_2298; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2301 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_2_6 : dataModule_io_maskOut_0_2_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2302 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_2_6 : _GEN_2301; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2303 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_2_6 : _GEN_2302; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2304 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_2_6 : _GEN_2303; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2305 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_2_6 : _GEN_2304; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2306 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_2_6 : _GEN_2305; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2307 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_2_6 : _GEN_2306; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2308 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_2_6 : _GEN_2307; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2309 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_2_6 : _GEN_2308; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2310 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_2_6 : _GEN_2309; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2311 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_2_6 : _GEN_2310; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2312 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_2_6 : _GEN_2311; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2313 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_2_6 : _GEN_2312; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2314 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_2_6 : _GEN_2313; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2315 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_2_6 : _GEN_2314; // @[Sbuffer.scala 704:{64,64}]
  wire [7:0] io_dcache_req_bits_mask_lo_hi_lo = {_GEN_2299,_GEN_2315,_GEN_2267,_GEN_2283,_GEN_2235,_GEN_2251,_GEN_2203,
    _GEN_2219}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2317 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_1 : dataModule_io_maskOut_0_3_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2318 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_1 : _GEN_2317; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2319 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_1 : _GEN_2318; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2320 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_1 : _GEN_2319; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2321 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_1 : _GEN_2320; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2322 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_1 : _GEN_2321; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2323 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_1 : _GEN_2322; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2324 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_1 : _GEN_2323; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2325 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_1 : _GEN_2324; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2326 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_1 : _GEN_2325; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2327 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_1 : _GEN_2326; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2328 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_1 : _GEN_2327; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2329 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_1 : _GEN_2328; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2330 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_1 : _GEN_2329; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2331 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_1 : _GEN_2330; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2333 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_0 : dataModule_io_maskOut_0_3_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2334 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_0 : _GEN_2333; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2335 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_0 : _GEN_2334; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2336 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_0 : _GEN_2335; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2337 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_0 : _GEN_2336; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2338 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_0 : _GEN_2337; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2339 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_0 : _GEN_2338; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2340 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_0 : _GEN_2339; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2341 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_0 : _GEN_2340; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2342 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_0 : _GEN_2341; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2343 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_0 : _GEN_2342; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2344 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_0 : _GEN_2343; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2345 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_0 : _GEN_2344; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2346 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_0 : _GEN_2345; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2347 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_0 : _GEN_2346; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2349 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_3 : dataModule_io_maskOut_0_3_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2350 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_3 : _GEN_2349; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2351 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_3 : _GEN_2350; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2352 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_3 : _GEN_2351; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2353 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_3 : _GEN_2352; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2354 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_3 : _GEN_2353; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2355 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_3 : _GEN_2354; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2356 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_3 : _GEN_2355; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2357 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_3 : _GEN_2356; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2358 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_3 : _GEN_2357; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2359 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_3 : _GEN_2358; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2360 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_3 : _GEN_2359; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2361 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_3 : _GEN_2360; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2362 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_3 : _GEN_2361; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2363 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_3 : _GEN_2362; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2365 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_2 : dataModule_io_maskOut_0_3_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2366 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_2 : _GEN_2365; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2367 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_2 : _GEN_2366; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2368 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_2 : _GEN_2367; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2369 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_2 : _GEN_2368; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2370 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_2 : _GEN_2369; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2371 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_2 : _GEN_2370; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2372 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_2 : _GEN_2371; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2373 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_2 : _GEN_2372; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2374 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_2 : _GEN_2373; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2375 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_2 : _GEN_2374; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2376 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_2 : _GEN_2375; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2377 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_2 : _GEN_2376; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2378 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_2 : _GEN_2377; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2379 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_2 : _GEN_2378; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2381 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_5 : dataModule_io_maskOut_0_3_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2382 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_5 : _GEN_2381; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2383 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_5 : _GEN_2382; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2384 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_5 : _GEN_2383; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2385 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_5 : _GEN_2384; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2386 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_5 : _GEN_2385; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2387 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_5 : _GEN_2386; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2388 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_5 : _GEN_2387; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2389 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_5 : _GEN_2388; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2390 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_5 : _GEN_2389; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2391 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_5 : _GEN_2390; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2392 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_5 : _GEN_2391; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2393 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_5 : _GEN_2392; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2394 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_5 : _GEN_2393; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2395 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_5 : _GEN_2394; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2397 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_4 : dataModule_io_maskOut_0_3_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2398 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_4 : _GEN_2397; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2399 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_4 : _GEN_2398; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2400 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_4 : _GEN_2399; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2401 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_4 : _GEN_2400; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2402 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_4 : _GEN_2401; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2403 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_4 : _GEN_2402; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2404 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_4 : _GEN_2403; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2405 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_4 : _GEN_2404; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2406 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_4 : _GEN_2405; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2407 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_4 : _GEN_2406; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2408 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_4 : _GEN_2407; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2409 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_4 : _GEN_2408; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2410 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_4 : _GEN_2409; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2411 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_4 : _GEN_2410; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2413 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_7 : dataModule_io_maskOut_0_3_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2414 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_7 : _GEN_2413; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2415 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_7 : _GEN_2414; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2416 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_7 : _GEN_2415; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2417 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_7 : _GEN_2416; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2418 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_7 : _GEN_2417; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2419 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_7 : _GEN_2418; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2420 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_7 : _GEN_2419; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2421 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_7 : _GEN_2420; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2422 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_7 : _GEN_2421; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2423 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_7 : _GEN_2422; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2424 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_7 : _GEN_2423; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2425 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_7 : _GEN_2424; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2426 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_7 : _GEN_2425; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2427 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_7 : _GEN_2426; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2429 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_3_6 : dataModule_io_maskOut_0_3_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2430 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_3_6 : _GEN_2429; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2431 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_3_6 : _GEN_2430; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2432 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_3_6 : _GEN_2431; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2433 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_3_6 : _GEN_2432; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2434 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_3_6 : _GEN_2433; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2435 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_3_6 : _GEN_2434; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2436 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_3_6 : _GEN_2435; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2437 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_3_6 : _GEN_2436; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2438 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_3_6 : _GEN_2437; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2439 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_3_6 : _GEN_2438; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2440 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_3_6 : _GEN_2439; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2441 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_3_6 : _GEN_2440; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2442 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_3_6 : _GEN_2441; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2443 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_3_6 : _GEN_2442; // @[Sbuffer.scala 704:{64,64}]
  wire [31:0] io_dcache_req_bits_mask_lo = {_GEN_2427,_GEN_2443,_GEN_2395,_GEN_2411,_GEN_2363,_GEN_2379,_GEN_2331,
    _GEN_2347,io_dcache_req_bits_mask_lo_hi_lo,io_dcache_req_bits_mask_lo_lo}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2445 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_1 : dataModule_io_maskOut_0_4_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2446 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_1 : _GEN_2445; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2447 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_1 : _GEN_2446; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2448 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_1 : _GEN_2447; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2449 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_1 : _GEN_2448; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2450 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_1 : _GEN_2449; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2451 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_1 : _GEN_2450; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2452 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_1 : _GEN_2451; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2453 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_1 : _GEN_2452; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2454 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_1 : _GEN_2453; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2455 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_1 : _GEN_2454; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2456 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_1 : _GEN_2455; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2457 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_1 : _GEN_2456; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2458 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_1 : _GEN_2457; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2459 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_1 : _GEN_2458; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2461 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_0 : dataModule_io_maskOut_0_4_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2462 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_0 : _GEN_2461; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2463 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_0 : _GEN_2462; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2464 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_0 : _GEN_2463; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2465 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_0 : _GEN_2464; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2466 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_0 : _GEN_2465; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2467 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_0 : _GEN_2466; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2468 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_0 : _GEN_2467; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2469 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_0 : _GEN_2468; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2470 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_0 : _GEN_2469; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2471 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_0 : _GEN_2470; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2472 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_0 : _GEN_2471; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2473 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_0 : _GEN_2472; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2474 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_0 : _GEN_2473; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2475 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_0 : _GEN_2474; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2477 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_3 : dataModule_io_maskOut_0_4_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2478 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_3 : _GEN_2477; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2479 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_3 : _GEN_2478; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2480 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_3 : _GEN_2479; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2481 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_3 : _GEN_2480; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2482 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_3 : _GEN_2481; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2483 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_3 : _GEN_2482; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2484 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_3 : _GEN_2483; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2485 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_3 : _GEN_2484; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2486 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_3 : _GEN_2485; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2487 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_3 : _GEN_2486; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2488 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_3 : _GEN_2487; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2489 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_3 : _GEN_2488; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2490 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_3 : _GEN_2489; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2491 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_3 : _GEN_2490; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2493 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_2 : dataModule_io_maskOut_0_4_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2494 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_2 : _GEN_2493; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2495 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_2 : _GEN_2494; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2496 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_2 : _GEN_2495; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2497 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_2 : _GEN_2496; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2498 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_2 : _GEN_2497; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2499 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_2 : _GEN_2498; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2500 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_2 : _GEN_2499; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2501 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_2 : _GEN_2500; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2502 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_2 : _GEN_2501; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2503 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_2 : _GEN_2502; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2504 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_2 : _GEN_2503; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2505 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_2 : _GEN_2504; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2506 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_2 : _GEN_2505; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2507 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_2 : _GEN_2506; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2509 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_5 : dataModule_io_maskOut_0_4_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2510 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_5 : _GEN_2509; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2511 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_5 : _GEN_2510; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2512 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_5 : _GEN_2511; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2513 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_5 : _GEN_2512; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2514 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_5 : _GEN_2513; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2515 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_5 : _GEN_2514; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2516 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_5 : _GEN_2515; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2517 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_5 : _GEN_2516; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2518 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_5 : _GEN_2517; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2519 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_5 : _GEN_2518; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2520 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_5 : _GEN_2519; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2521 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_5 : _GEN_2520; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2522 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_5 : _GEN_2521; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2523 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_5 : _GEN_2522; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2525 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_4 : dataModule_io_maskOut_0_4_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2526 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_4 : _GEN_2525; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2527 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_4 : _GEN_2526; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2528 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_4 : _GEN_2527; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2529 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_4 : _GEN_2528; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2530 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_4 : _GEN_2529; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2531 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_4 : _GEN_2530; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2532 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_4 : _GEN_2531; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2533 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_4 : _GEN_2532; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2534 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_4 : _GEN_2533; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2535 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_4 : _GEN_2534; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2536 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_4 : _GEN_2535; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2537 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_4 : _GEN_2536; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2538 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_4 : _GEN_2537; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2539 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_4 : _GEN_2538; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2541 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_7 : dataModule_io_maskOut_0_4_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2542 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_7 : _GEN_2541; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2543 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_7 : _GEN_2542; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2544 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_7 : _GEN_2543; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2545 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_7 : _GEN_2544; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2546 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_7 : _GEN_2545; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2547 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_7 : _GEN_2546; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2548 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_7 : _GEN_2547; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2549 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_7 : _GEN_2548; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2550 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_7 : _GEN_2549; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2551 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_7 : _GEN_2550; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2552 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_7 : _GEN_2551; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2553 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_7 : _GEN_2552; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2554 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_7 : _GEN_2553; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2555 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_7 : _GEN_2554; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2557 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_4_6 : dataModule_io_maskOut_0_4_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2558 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_4_6 : _GEN_2557; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2559 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_4_6 : _GEN_2558; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2560 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_4_6 : _GEN_2559; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2561 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_4_6 : _GEN_2560; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2562 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_4_6 : _GEN_2561; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2563 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_4_6 : _GEN_2562; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2564 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_4_6 : _GEN_2563; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2565 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_4_6 : _GEN_2564; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2566 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_4_6 : _GEN_2565; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2567 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_4_6 : _GEN_2566; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2568 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_4_6 : _GEN_2567; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2569 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_4_6 : _GEN_2568; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2570 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_4_6 : _GEN_2569; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2571 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_4_6 : _GEN_2570; // @[Sbuffer.scala 704:{64,64}]
  wire [7:0] io_dcache_req_bits_mask_hi_lo_lo = {_GEN_2555,_GEN_2571,_GEN_2523,_GEN_2539,_GEN_2491,_GEN_2507,_GEN_2459,
    _GEN_2475}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2573 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_1 : dataModule_io_maskOut_0_5_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2574 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_1 : _GEN_2573; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2575 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_1 : _GEN_2574; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2576 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_1 : _GEN_2575; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2577 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_1 : _GEN_2576; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2578 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_1 : _GEN_2577; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2579 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_1 : _GEN_2578; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2580 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_1 : _GEN_2579; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2581 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_1 : _GEN_2580; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2582 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_1 : _GEN_2581; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2583 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_1 : _GEN_2582; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2584 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_1 : _GEN_2583; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2585 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_1 : _GEN_2584; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2586 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_1 : _GEN_2585; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2587 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_1 : _GEN_2586; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2589 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_0 : dataModule_io_maskOut_0_5_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2590 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_0 : _GEN_2589; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2591 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_0 : _GEN_2590; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2592 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_0 : _GEN_2591; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2593 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_0 : _GEN_2592; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2594 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_0 : _GEN_2593; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2595 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_0 : _GEN_2594; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2596 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_0 : _GEN_2595; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2597 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_0 : _GEN_2596; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2598 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_0 : _GEN_2597; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2599 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_0 : _GEN_2598; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2600 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_0 : _GEN_2599; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2601 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_0 : _GEN_2600; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2602 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_0 : _GEN_2601; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2603 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_0 : _GEN_2602; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2605 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_3 : dataModule_io_maskOut_0_5_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2606 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_3 : _GEN_2605; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2607 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_3 : _GEN_2606; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2608 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_3 : _GEN_2607; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2609 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_3 : _GEN_2608; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2610 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_3 : _GEN_2609; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2611 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_3 : _GEN_2610; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2612 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_3 : _GEN_2611; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2613 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_3 : _GEN_2612; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2614 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_3 : _GEN_2613; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2615 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_3 : _GEN_2614; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2616 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_3 : _GEN_2615; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2617 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_3 : _GEN_2616; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2618 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_3 : _GEN_2617; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2619 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_3 : _GEN_2618; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2621 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_2 : dataModule_io_maskOut_0_5_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2622 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_2 : _GEN_2621; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2623 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_2 : _GEN_2622; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2624 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_2 : _GEN_2623; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2625 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_2 : _GEN_2624; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2626 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_2 : _GEN_2625; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2627 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_2 : _GEN_2626; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2628 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_2 : _GEN_2627; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2629 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_2 : _GEN_2628; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2630 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_2 : _GEN_2629; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2631 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_2 : _GEN_2630; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2632 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_2 : _GEN_2631; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2633 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_2 : _GEN_2632; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2634 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_2 : _GEN_2633; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2635 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_2 : _GEN_2634; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2637 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_5 : dataModule_io_maskOut_0_5_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2638 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_5 : _GEN_2637; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2639 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_5 : _GEN_2638; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2640 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_5 : _GEN_2639; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2641 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_5 : _GEN_2640; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2642 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_5 : _GEN_2641; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2643 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_5 : _GEN_2642; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2644 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_5 : _GEN_2643; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2645 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_5 : _GEN_2644; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2646 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_5 : _GEN_2645; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2647 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_5 : _GEN_2646; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2648 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_5 : _GEN_2647; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2649 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_5 : _GEN_2648; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2650 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_5 : _GEN_2649; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2651 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_5 : _GEN_2650; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2653 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_4 : dataModule_io_maskOut_0_5_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2654 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_4 : _GEN_2653; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2655 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_4 : _GEN_2654; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2656 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_4 : _GEN_2655; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2657 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_4 : _GEN_2656; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2658 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_4 : _GEN_2657; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2659 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_4 : _GEN_2658; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2660 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_4 : _GEN_2659; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2661 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_4 : _GEN_2660; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2662 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_4 : _GEN_2661; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2663 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_4 : _GEN_2662; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2664 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_4 : _GEN_2663; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2665 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_4 : _GEN_2664; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2666 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_4 : _GEN_2665; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2667 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_4 : _GEN_2666; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2669 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_7 : dataModule_io_maskOut_0_5_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2670 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_7 : _GEN_2669; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2671 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_7 : _GEN_2670; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2672 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_7 : _GEN_2671; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2673 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_7 : _GEN_2672; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2674 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_7 : _GEN_2673; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2675 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_7 : _GEN_2674; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2676 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_7 : _GEN_2675; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2677 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_7 : _GEN_2676; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2678 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_7 : _GEN_2677; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2679 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_7 : _GEN_2678; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2680 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_7 : _GEN_2679; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2681 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_7 : _GEN_2680; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2682 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_7 : _GEN_2681; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2683 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_7 : _GEN_2682; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2685 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_5_6 : dataModule_io_maskOut_0_5_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2686 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_5_6 : _GEN_2685; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2687 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_5_6 : _GEN_2686; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2688 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_5_6 : _GEN_2687; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2689 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_5_6 : _GEN_2688; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2690 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_5_6 : _GEN_2689; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2691 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_5_6 : _GEN_2690; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2692 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_5_6 : _GEN_2691; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2693 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_5_6 : _GEN_2692; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2694 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_5_6 : _GEN_2693; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2695 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_5_6 : _GEN_2694; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2696 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_5_6 : _GEN_2695; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2697 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_5_6 : _GEN_2696; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2698 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_5_6 : _GEN_2697; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2699 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_5_6 : _GEN_2698; // @[Sbuffer.scala 704:{64,64}]
  wire [15:0] io_dcache_req_bits_mask_hi_lo = {_GEN_2683,_GEN_2699,_GEN_2651,_GEN_2667,_GEN_2619,_GEN_2635,_GEN_2587,
    _GEN_2603,io_dcache_req_bits_mask_hi_lo_lo}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2701 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_1 : dataModule_io_maskOut_0_6_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2702 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_1 : _GEN_2701; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2703 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_1 : _GEN_2702; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2704 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_1 : _GEN_2703; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2705 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_1 : _GEN_2704; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2706 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_1 : _GEN_2705; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2707 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_1 : _GEN_2706; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2708 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_1 : _GEN_2707; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2709 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_1 : _GEN_2708; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2710 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_1 : _GEN_2709; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2711 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_1 : _GEN_2710; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2712 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_1 : _GEN_2711; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2713 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_1 : _GEN_2712; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2714 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_1 : _GEN_2713; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2715 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_1 : _GEN_2714; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2717 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_0 : dataModule_io_maskOut_0_6_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2718 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_0 : _GEN_2717; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2719 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_0 : _GEN_2718; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2720 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_0 : _GEN_2719; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2721 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_0 : _GEN_2720; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2722 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_0 : _GEN_2721; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2723 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_0 : _GEN_2722; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2724 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_0 : _GEN_2723; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2725 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_0 : _GEN_2724; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2726 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_0 : _GEN_2725; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2727 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_0 : _GEN_2726; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2728 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_0 : _GEN_2727; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2729 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_0 : _GEN_2728; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2730 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_0 : _GEN_2729; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2731 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_0 : _GEN_2730; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2733 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_3 : dataModule_io_maskOut_0_6_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2734 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_3 : _GEN_2733; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2735 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_3 : _GEN_2734; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2736 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_3 : _GEN_2735; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2737 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_3 : _GEN_2736; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2738 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_3 : _GEN_2737; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2739 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_3 : _GEN_2738; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2740 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_3 : _GEN_2739; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2741 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_3 : _GEN_2740; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2742 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_3 : _GEN_2741; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2743 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_3 : _GEN_2742; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2744 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_3 : _GEN_2743; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2745 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_3 : _GEN_2744; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2746 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_3 : _GEN_2745; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2747 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_3 : _GEN_2746; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2749 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_2 : dataModule_io_maskOut_0_6_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2750 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_2 : _GEN_2749; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2751 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_2 : _GEN_2750; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2752 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_2 : _GEN_2751; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2753 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_2 : _GEN_2752; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2754 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_2 : _GEN_2753; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2755 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_2 : _GEN_2754; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2756 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_2 : _GEN_2755; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2757 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_2 : _GEN_2756; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2758 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_2 : _GEN_2757; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2759 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_2 : _GEN_2758; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2760 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_2 : _GEN_2759; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2761 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_2 : _GEN_2760; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2762 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_2 : _GEN_2761; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2763 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_2 : _GEN_2762; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2765 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_5 : dataModule_io_maskOut_0_6_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2766 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_5 : _GEN_2765; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2767 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_5 : _GEN_2766; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2768 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_5 : _GEN_2767; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2769 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_5 : _GEN_2768; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2770 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_5 : _GEN_2769; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2771 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_5 : _GEN_2770; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2772 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_5 : _GEN_2771; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2773 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_5 : _GEN_2772; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2774 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_5 : _GEN_2773; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2775 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_5 : _GEN_2774; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2776 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_5 : _GEN_2775; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2777 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_5 : _GEN_2776; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2778 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_5 : _GEN_2777; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2779 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_5 : _GEN_2778; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2781 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_4 : dataModule_io_maskOut_0_6_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2782 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_4 : _GEN_2781; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2783 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_4 : _GEN_2782; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2784 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_4 : _GEN_2783; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2785 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_4 : _GEN_2784; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2786 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_4 : _GEN_2785; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2787 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_4 : _GEN_2786; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2788 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_4 : _GEN_2787; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2789 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_4 : _GEN_2788; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2790 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_4 : _GEN_2789; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2791 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_4 : _GEN_2790; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2792 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_4 : _GEN_2791; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2793 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_4 : _GEN_2792; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2794 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_4 : _GEN_2793; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2795 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_4 : _GEN_2794; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2797 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_7 : dataModule_io_maskOut_0_6_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2798 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_7 : _GEN_2797; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2799 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_7 : _GEN_2798; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2800 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_7 : _GEN_2799; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2801 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_7 : _GEN_2800; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2802 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_7 : _GEN_2801; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2803 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_7 : _GEN_2802; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2804 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_7 : _GEN_2803; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2805 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_7 : _GEN_2804; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2806 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_7 : _GEN_2805; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2807 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_7 : _GEN_2806; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2808 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_7 : _GEN_2807; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2809 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_7 : _GEN_2808; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2810 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_7 : _GEN_2809; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2811 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_7 : _GEN_2810; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2813 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_6_6 : dataModule_io_maskOut_0_6_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2814 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_6_6 : _GEN_2813; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2815 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_6_6 : _GEN_2814; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2816 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_6_6 : _GEN_2815; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2817 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_6_6 : _GEN_2816; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2818 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_6_6 : _GEN_2817; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2819 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_6_6 : _GEN_2818; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2820 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_6_6 : _GEN_2819; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2821 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_6_6 : _GEN_2820; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2822 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_6_6 : _GEN_2821; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2823 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_6_6 : _GEN_2822; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2824 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_6_6 : _GEN_2823; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2825 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_6_6 : _GEN_2824; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2826 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_6_6 : _GEN_2825; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2827 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_6_6 : _GEN_2826; // @[Sbuffer.scala 704:{64,64}]
  wire [7:0] io_dcache_req_bits_mask_hi_hi_lo = {_GEN_2811,_GEN_2827,_GEN_2779,_GEN_2795,_GEN_2747,_GEN_2763,_GEN_2715,
    _GEN_2731}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2829 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_1 : dataModule_io_maskOut_0_7_1; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2830 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_1 : _GEN_2829; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2831 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_1 : _GEN_2830; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2832 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_1 : _GEN_2831; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2833 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_1 : _GEN_2832; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2834 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_1 : _GEN_2833; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2835 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_1 : _GEN_2834; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2836 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_1 : _GEN_2835; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2837 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_1 : _GEN_2836; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2838 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_1 : _GEN_2837; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2839 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_1 : _GEN_2838; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2840 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_1 : _GEN_2839; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2841 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_1 : _GEN_2840; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2842 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_1 : _GEN_2841; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2843 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_1 : _GEN_2842; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2845 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_0 : dataModule_io_maskOut_0_7_0; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2846 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_0 : _GEN_2845; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2847 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_0 : _GEN_2846; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2848 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_0 : _GEN_2847; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2849 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_0 : _GEN_2848; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2850 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_0 : _GEN_2849; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2851 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_0 : _GEN_2850; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2852 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_0 : _GEN_2851; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2853 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_0 : _GEN_2852; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2854 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_0 : _GEN_2853; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2855 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_0 : _GEN_2854; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2856 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_0 : _GEN_2855; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2857 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_0 : _GEN_2856; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2858 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_0 : _GEN_2857; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2859 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_0 : _GEN_2858; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2861 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_3 : dataModule_io_maskOut_0_7_3; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2862 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_3 : _GEN_2861; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2863 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_3 : _GEN_2862; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2864 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_3 : _GEN_2863; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2865 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_3 : _GEN_2864; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2866 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_3 : _GEN_2865; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2867 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_3 : _GEN_2866; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2868 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_3 : _GEN_2867; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2869 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_3 : _GEN_2868; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2870 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_3 : _GEN_2869; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2871 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_3 : _GEN_2870; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2872 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_3 : _GEN_2871; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2873 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_3 : _GEN_2872; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2874 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_3 : _GEN_2873; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2875 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_3 : _GEN_2874; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2877 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_2 : dataModule_io_maskOut_0_7_2; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2878 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_2 : _GEN_2877; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2879 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_2 : _GEN_2878; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2880 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_2 : _GEN_2879; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2881 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_2 : _GEN_2880; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2882 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_2 : _GEN_2881; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2883 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_2 : _GEN_2882; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2884 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_2 : _GEN_2883; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2885 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_2 : _GEN_2884; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2886 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_2 : _GEN_2885; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2887 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_2 : _GEN_2886; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2888 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_2 : _GEN_2887; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2889 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_2 : _GEN_2888; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2890 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_2 : _GEN_2889; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2891 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_2 : _GEN_2890; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2893 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_5 : dataModule_io_maskOut_0_7_5; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2894 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_5 : _GEN_2893; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2895 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_5 : _GEN_2894; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2896 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_5 : _GEN_2895; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2897 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_5 : _GEN_2896; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2898 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_5 : _GEN_2897; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2899 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_5 : _GEN_2898; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2900 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_5 : _GEN_2899; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2901 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_5 : _GEN_2900; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2902 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_5 : _GEN_2901; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2903 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_5 : _GEN_2902; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2904 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_5 : _GEN_2903; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2905 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_5 : _GEN_2904; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2906 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_5 : _GEN_2905; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2907 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_5 : _GEN_2906; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2909 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_4 : dataModule_io_maskOut_0_7_4; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2910 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_4 : _GEN_2909; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2911 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_4 : _GEN_2910; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2912 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_4 : _GEN_2911; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2913 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_4 : _GEN_2912; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2914 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_4 : _GEN_2913; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2915 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_4 : _GEN_2914; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2916 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_4 : _GEN_2915; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2917 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_4 : _GEN_2916; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2918 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_4 : _GEN_2917; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2919 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_4 : _GEN_2918; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2920 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_4 : _GEN_2919; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2921 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_4 : _GEN_2920; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2922 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_4 : _GEN_2921; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2923 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_4 : _GEN_2922; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2925 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_7 : dataModule_io_maskOut_0_7_7; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2926 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_7 : _GEN_2925; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2927 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_7 : _GEN_2926; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2928 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_7 : _GEN_2927; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2929 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_7 : _GEN_2928; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2930 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_7 : _GEN_2929; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2931 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_7 : _GEN_2930; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2932 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_7 : _GEN_2931; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2933 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_7 : _GEN_2932; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2934 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_7 : _GEN_2933; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2935 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_7 : _GEN_2934; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2936 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_7 : _GEN_2935; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2937 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_7 : _GEN_2936; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2938 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_7 : _GEN_2937; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2939 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_7 : _GEN_2938; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2941 = 4'h1 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_1_7_6 : dataModule_io_maskOut_0_7_6; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2942 = 4'h2 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_2_7_6 : _GEN_2941; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2943 = 4'h3 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_3_7_6 : _GEN_2942; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2944 = 4'h4 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_4_7_6 : _GEN_2943; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2945 = 4'h5 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_5_7_6 : _GEN_2944; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2946 = 4'h6 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_6_7_6 : _GEN_2945; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2947 = 4'h7 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_7_7_6 : _GEN_2946; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2948 = 4'h8 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_8_7_6 : _GEN_2947; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2949 = 4'h9 == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_9_7_6 : _GEN_2948; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2950 = 4'ha == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_10_7_6 : _GEN_2949; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2951 = 4'hb == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_11_7_6 : _GEN_2950; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2952 = 4'hc == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_12_7_6 : _GEN_2951; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2953 = 4'hd == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_13_7_6 : _GEN_2952; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2954 = 4'he == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_14_7_6 : _GEN_2953; // @[Sbuffer.scala 704:{64,64}]
  wire  _GEN_2955 = 4'hf == sbuffer_out_s1_evictionIdx ? dataModule_io_maskOut_15_7_6 : _GEN_2954; // @[Sbuffer.scala 704:{64,64}]
  wire [31:0] io_dcache_req_bits_mask_hi = {_GEN_2939,_GEN_2955,_GEN_2907,_GEN_2923,_GEN_2875,_GEN_2891,_GEN_2843,
    _GEN_2859,io_dcache_req_bits_mask_hi_hi_lo,io_dcache_req_bits_mask_hi_lo}; // @[Sbuffer.scala 704:64]
  wire  _GEN_2956 = 4'h0 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_825; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2957 = 4'h1 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_826; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2958 = 4'h2 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_827; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2959 = 4'h3 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_828; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2960 = 4'h4 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_829; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2961 = 4'h5 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_830; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2962 = 4'h6 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_831; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2963 = 4'h7 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_832; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2964 = 4'h8 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_833; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2965 = 4'h9 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_834; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2966 = 4'ha == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_835; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2967 = 4'hb == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_836; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2968 = 4'hc == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_837; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2969 = 4'hd == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_838; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2970 = 4'he == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_839; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2971 = 4'hf == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_840; // @[Sbuffer.scala 727:{47,47}]
  wire  _GEN_2972 = 4'h0 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_634; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2973 = 4'h1 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_639; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2974 = 4'h2 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_644; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2975 = 4'h3 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_649; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2976 = 4'h4 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_654; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2977 = 4'h5 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_659; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2978 = 4'h6 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_664; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2979 = 4'h7 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_669; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2980 = 4'h8 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_674; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2981 = 4'h9 == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_679; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2982 = 4'ha == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_684; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2983 = 4'hb == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_689; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2984 = 4'hc == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_694; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2985 = 4'hd == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_699; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2986 = 4'he == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_704; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_2987 = 4'hf == io_dcache_main_pipe_hit_resp_bits_id[3:0] ? 1'h0 : _GEN_709; // @[Sbuffer.scala 728:{44,44}]
  wire  _GEN_3004 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2956 : _GEN_825; // @[Sbuffer.scala 726:24]
  wire  _GEN_3005 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2957 : _GEN_826; // @[Sbuffer.scala 726:24]
  wire  _GEN_3006 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2958 : _GEN_827; // @[Sbuffer.scala 726:24]
  wire  _GEN_3007 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2959 : _GEN_828; // @[Sbuffer.scala 726:24]
  wire  _GEN_3008 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2960 : _GEN_829; // @[Sbuffer.scala 726:24]
  wire  _GEN_3009 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2961 : _GEN_830; // @[Sbuffer.scala 726:24]
  wire  _GEN_3010 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2962 : _GEN_831; // @[Sbuffer.scala 726:24]
  wire  _GEN_3011 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2963 : _GEN_832; // @[Sbuffer.scala 726:24]
  wire  _GEN_3012 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2964 : _GEN_833; // @[Sbuffer.scala 726:24]
  wire  _GEN_3013 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2965 : _GEN_834; // @[Sbuffer.scala 726:24]
  wire  _GEN_3014 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2966 : _GEN_835; // @[Sbuffer.scala 726:24]
  wire  _GEN_3015 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2967 : _GEN_836; // @[Sbuffer.scala 726:24]
  wire  _GEN_3016 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2968 : _GEN_837; // @[Sbuffer.scala 726:24]
  wire  _GEN_3017 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2969 : _GEN_838; // @[Sbuffer.scala 726:24]
  wire  _GEN_3018 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2970 : _GEN_839; // @[Sbuffer.scala 726:24]
  wire  _GEN_3019 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2971 : _GEN_840; // @[Sbuffer.scala 726:24]
  wire  _GEN_3020 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2972 : _GEN_634; // @[Sbuffer.scala 726:24]
  wire  _GEN_3021 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2973 : _GEN_639; // @[Sbuffer.scala 726:24]
  wire  _GEN_3022 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2974 : _GEN_644; // @[Sbuffer.scala 726:24]
  wire  _GEN_3023 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2975 : _GEN_649; // @[Sbuffer.scala 726:24]
  wire  _GEN_3024 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2976 : _GEN_654; // @[Sbuffer.scala 726:24]
  wire  _GEN_3025 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2977 : _GEN_659; // @[Sbuffer.scala 726:24]
  wire  _GEN_3026 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2978 : _GEN_664; // @[Sbuffer.scala 726:24]
  wire  _GEN_3027 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2979 : _GEN_669; // @[Sbuffer.scala 726:24]
  wire  _GEN_3028 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2980 : _GEN_674; // @[Sbuffer.scala 726:24]
  wire  _GEN_3029 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2981 : _GEN_679; // @[Sbuffer.scala 726:24]
  wire  _GEN_3030 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2982 : _GEN_684; // @[Sbuffer.scala 726:24]
  wire  _GEN_3031 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2983 : _GEN_689; // @[Sbuffer.scala 726:24]
  wire  _GEN_3032 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2984 : _GEN_694; // @[Sbuffer.scala 726:24]
  wire  _GEN_3033 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2985 : _GEN_699; // @[Sbuffer.scala 726:24]
  wire  _GEN_3034 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2986 : _GEN_704; // @[Sbuffer.scala 726:24]
  wire  _GEN_3035 = io_dcache_main_pipe_hit_resp_valid ? _GEN_2987 : _GEN_709; // @[Sbuffer.scala 726:24]
  wire  _T_713 = stateVec_0_w_sameblock_inflight & stateVec_0_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG; // @[Sbuffer.scala 743:16]
  wire  _T_714 = _T_713 & REG; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_1; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_716 = 16'h1 << REG_1; // @[OneHot.scala 57:35]
  wire  _T_717 = waitInflightMask_0 == _T_716; // @[Sbuffer.scala 744:29]
  wire  _T_718 = _T_714 & _T_717; // @[Sbuffer.scala 743:30]
  wire  _T_719 = stateVec_1_w_sameblock_inflight & stateVec_1_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_2; // @[Sbuffer.scala 743:16]
  wire  _T_720 = _T_719 & REG_2; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_3; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_722 = 16'h1 << REG_3; // @[OneHot.scala 57:35]
  wire  _T_723 = waitInflightMask_1 == _T_722; // @[Sbuffer.scala 744:29]
  wire  _T_724 = _T_720 & _T_723; // @[Sbuffer.scala 743:30]
  wire  _T_725 = stateVec_2_w_sameblock_inflight & stateVec_2_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_4; // @[Sbuffer.scala 743:16]
  wire  _T_726 = _T_725 & REG_4; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_5; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_728 = 16'h1 << REG_5; // @[OneHot.scala 57:35]
  wire  _T_729 = waitInflightMask_2 == _T_728; // @[Sbuffer.scala 744:29]
  wire  _T_730 = _T_726 & _T_729; // @[Sbuffer.scala 743:30]
  wire  _T_731 = stateVec_3_w_sameblock_inflight & stateVec_3_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_6; // @[Sbuffer.scala 743:16]
  wire  _T_732 = _T_731 & REG_6; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_7; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_734 = 16'h1 << REG_7; // @[OneHot.scala 57:35]
  wire  _T_735 = waitInflightMask_3 == _T_734; // @[Sbuffer.scala 744:29]
  wire  _T_736 = _T_732 & _T_735; // @[Sbuffer.scala 743:30]
  wire  _T_737 = stateVec_4_w_sameblock_inflight & stateVec_4_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_8; // @[Sbuffer.scala 743:16]
  wire  _T_738 = _T_737 & REG_8; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_9; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_740 = 16'h1 << REG_9; // @[OneHot.scala 57:35]
  wire  _T_741 = waitInflightMask_4 == _T_740; // @[Sbuffer.scala 744:29]
  wire  _T_742 = _T_738 & _T_741; // @[Sbuffer.scala 743:30]
  wire  _T_743 = stateVec_5_w_sameblock_inflight & stateVec_5_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_10; // @[Sbuffer.scala 743:16]
  wire  _T_744 = _T_743 & REG_10; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_11; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_746 = 16'h1 << REG_11; // @[OneHot.scala 57:35]
  wire  _T_747 = waitInflightMask_5 == _T_746; // @[Sbuffer.scala 744:29]
  wire  _T_748 = _T_744 & _T_747; // @[Sbuffer.scala 743:30]
  wire  _T_749 = stateVec_6_w_sameblock_inflight & stateVec_6_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_12; // @[Sbuffer.scala 743:16]
  wire  _T_750 = _T_749 & REG_12; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_13; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_752 = 16'h1 << REG_13; // @[OneHot.scala 57:35]
  wire  _T_753 = waitInflightMask_6 == _T_752; // @[Sbuffer.scala 744:29]
  wire  _T_754 = _T_750 & _T_753; // @[Sbuffer.scala 743:30]
  wire  _T_755 = stateVec_7_w_sameblock_inflight & stateVec_7_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_14; // @[Sbuffer.scala 743:16]
  wire  _T_756 = _T_755 & REG_14; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_15; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_758 = 16'h1 << REG_15; // @[OneHot.scala 57:35]
  wire  _T_759 = waitInflightMask_7 == _T_758; // @[Sbuffer.scala 744:29]
  wire  _T_760 = _T_756 & _T_759; // @[Sbuffer.scala 743:30]
  wire  _T_761 = stateVec_8_w_sameblock_inflight & stateVec_8_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_16; // @[Sbuffer.scala 743:16]
  wire  _T_762 = _T_761 & REG_16; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_17; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_764 = 16'h1 << REG_17; // @[OneHot.scala 57:35]
  wire  _T_765 = waitInflightMask_8 == _T_764; // @[Sbuffer.scala 744:29]
  wire  _T_766 = _T_762 & _T_765; // @[Sbuffer.scala 743:30]
  wire  _T_767 = stateVec_9_w_sameblock_inflight & stateVec_9_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_18; // @[Sbuffer.scala 743:16]
  wire  _T_768 = _T_767 & REG_18; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_19; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_770 = 16'h1 << REG_19; // @[OneHot.scala 57:35]
  wire  _T_771 = waitInflightMask_9 == _T_770; // @[Sbuffer.scala 744:29]
  wire  _T_772 = _T_768 & _T_771; // @[Sbuffer.scala 743:30]
  wire  _T_773 = stateVec_10_w_sameblock_inflight & stateVec_10_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_20; // @[Sbuffer.scala 743:16]
  wire  _T_774 = _T_773 & REG_20; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_21; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_776 = 16'h1 << REG_21; // @[OneHot.scala 57:35]
  wire  _T_777 = waitInflightMask_10 == _T_776; // @[Sbuffer.scala 744:29]
  wire  _T_778 = _T_774 & _T_777; // @[Sbuffer.scala 743:30]
  wire  _T_779 = stateVec_11_w_sameblock_inflight & stateVec_11_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_22; // @[Sbuffer.scala 743:16]
  wire  _T_780 = _T_779 & REG_22; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_23; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_782 = 16'h1 << REG_23; // @[OneHot.scala 57:35]
  wire  _T_783 = waitInflightMask_11 == _T_782; // @[Sbuffer.scala 744:29]
  wire  _T_784 = _T_780 & _T_783; // @[Sbuffer.scala 743:30]
  wire  _T_785 = stateVec_12_w_sameblock_inflight & stateVec_12_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_24; // @[Sbuffer.scala 743:16]
  wire  _T_786 = _T_785 & REG_24; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_25; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_788 = 16'h1 << REG_25; // @[OneHot.scala 57:35]
  wire  _T_789 = waitInflightMask_12 == _T_788; // @[Sbuffer.scala 744:29]
  wire  _T_790 = _T_786 & _T_789; // @[Sbuffer.scala 743:30]
  wire  _T_791 = stateVec_13_w_sameblock_inflight & stateVec_13_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_26; // @[Sbuffer.scala 743:16]
  wire  _T_792 = _T_791 & REG_26; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_27; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_794 = 16'h1 << REG_27; // @[OneHot.scala 57:35]
  wire  _T_795 = waitInflightMask_13 == _T_794; // @[Sbuffer.scala 744:29]
  wire  _T_796 = _T_792 & _T_795; // @[Sbuffer.scala 743:30]
  wire  _T_797 = stateVec_14_w_sameblock_inflight & stateVec_14_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_28; // @[Sbuffer.scala 743:16]
  wire  _T_798 = _T_797 & REG_28; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_29; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_800 = 16'h1 << REG_29; // @[OneHot.scala 57:35]
  wire  _T_801 = waitInflightMask_14 == _T_800; // @[Sbuffer.scala 744:29]
  wire  _T_802 = _T_798 & _T_801; // @[Sbuffer.scala 743:30]
  wire  _T_803 = stateVec_15_w_sameblock_inflight & stateVec_15_state_valid; // @[Sbuffer.scala 741:42]
  reg  REG_30; // @[Sbuffer.scala 743:16]
  wire  _T_804 = _T_803 & REG_30; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_31; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_806 = 16'h1 << REG_31; // @[OneHot.scala 57:35]
  wire  _T_807 = waitInflightMask_15 == _T_806; // @[Sbuffer.scala 744:29]
  wire  _T_808 = _T_804 & _T_807; // @[Sbuffer.scala 743:30]
  reg  REG_32; // @[Sbuffer.scala 743:16]
  wire  _T_825 = _T_713 & REG_32; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_33; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_827 = 16'h1 << REG_33; // @[OneHot.scala 57:35]
  wire  _T_828 = waitInflightMask_0 == _T_827; // @[Sbuffer.scala 744:29]
  wire  _T_829 = _T_825 & _T_828; // @[Sbuffer.scala 743:30]
  reg  REG_34; // @[Sbuffer.scala 743:16]
  wire  _T_831 = _T_719 & REG_34; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_35; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_833 = 16'h1 << REG_35; // @[OneHot.scala 57:35]
  wire  _T_834 = waitInflightMask_1 == _T_833; // @[Sbuffer.scala 744:29]
  wire  _T_835 = _T_831 & _T_834; // @[Sbuffer.scala 743:30]
  reg  REG_36; // @[Sbuffer.scala 743:16]
  wire  _T_837 = _T_725 & REG_36; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_37; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_839 = 16'h1 << REG_37; // @[OneHot.scala 57:35]
  wire  _T_840 = waitInflightMask_2 == _T_839; // @[Sbuffer.scala 744:29]
  wire  _T_841 = _T_837 & _T_840; // @[Sbuffer.scala 743:30]
  reg  REG_38; // @[Sbuffer.scala 743:16]
  wire  _T_843 = _T_731 & REG_38; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_39; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_845 = 16'h1 << REG_39; // @[OneHot.scala 57:35]
  wire  _T_846 = waitInflightMask_3 == _T_845; // @[Sbuffer.scala 744:29]
  wire  _T_847 = _T_843 & _T_846; // @[Sbuffer.scala 743:30]
  reg  REG_40; // @[Sbuffer.scala 743:16]
  wire  _T_849 = _T_737 & REG_40; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_41; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_851 = 16'h1 << REG_41; // @[OneHot.scala 57:35]
  wire  _T_852 = waitInflightMask_4 == _T_851; // @[Sbuffer.scala 744:29]
  wire  _T_853 = _T_849 & _T_852; // @[Sbuffer.scala 743:30]
  reg  REG_42; // @[Sbuffer.scala 743:16]
  wire  _T_855 = _T_743 & REG_42; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_43; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_857 = 16'h1 << REG_43; // @[OneHot.scala 57:35]
  wire  _T_858 = waitInflightMask_5 == _T_857; // @[Sbuffer.scala 744:29]
  wire  _T_859 = _T_855 & _T_858; // @[Sbuffer.scala 743:30]
  reg  REG_44; // @[Sbuffer.scala 743:16]
  wire  _T_861 = _T_749 & REG_44; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_45; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_863 = 16'h1 << REG_45; // @[OneHot.scala 57:35]
  wire  _T_864 = waitInflightMask_6 == _T_863; // @[Sbuffer.scala 744:29]
  wire  _T_865 = _T_861 & _T_864; // @[Sbuffer.scala 743:30]
  reg  REG_46; // @[Sbuffer.scala 743:16]
  wire  _T_867 = _T_755 & REG_46; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_47; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_869 = 16'h1 << REG_47; // @[OneHot.scala 57:35]
  wire  _T_870 = waitInflightMask_7 == _T_869; // @[Sbuffer.scala 744:29]
  wire  _T_871 = _T_867 & _T_870; // @[Sbuffer.scala 743:30]
  reg  REG_48; // @[Sbuffer.scala 743:16]
  wire  _T_873 = _T_761 & REG_48; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_49; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_875 = 16'h1 << REG_49; // @[OneHot.scala 57:35]
  wire  _T_876 = waitInflightMask_8 == _T_875; // @[Sbuffer.scala 744:29]
  wire  _T_877 = _T_873 & _T_876; // @[Sbuffer.scala 743:30]
  reg  REG_50; // @[Sbuffer.scala 743:16]
  wire  _T_879 = _T_767 & REG_50; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_51; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_881 = 16'h1 << REG_51; // @[OneHot.scala 57:35]
  wire  _T_882 = waitInflightMask_9 == _T_881; // @[Sbuffer.scala 744:29]
  wire  _T_883 = _T_879 & _T_882; // @[Sbuffer.scala 743:30]
  reg  REG_52; // @[Sbuffer.scala 743:16]
  wire  _T_885 = _T_773 & REG_52; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_53; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_887 = 16'h1 << REG_53; // @[OneHot.scala 57:35]
  wire  _T_888 = waitInflightMask_10 == _T_887; // @[Sbuffer.scala 744:29]
  wire  _T_889 = _T_885 & _T_888; // @[Sbuffer.scala 743:30]
  reg  REG_54; // @[Sbuffer.scala 743:16]
  wire  _T_891 = _T_779 & REG_54; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_55; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_893 = 16'h1 << REG_55; // @[OneHot.scala 57:35]
  wire  _T_894 = waitInflightMask_11 == _T_893; // @[Sbuffer.scala 744:29]
  wire  _T_895 = _T_891 & _T_894; // @[Sbuffer.scala 743:30]
  reg  REG_56; // @[Sbuffer.scala 743:16]
  wire  _T_897 = _T_785 & REG_56; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_57; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_899 = 16'h1 << REG_57; // @[OneHot.scala 57:35]
  wire  _T_900 = waitInflightMask_12 == _T_899; // @[Sbuffer.scala 744:29]
  wire  _T_901 = _T_897 & _T_900; // @[Sbuffer.scala 743:30]
  reg  REG_58; // @[Sbuffer.scala 743:16]
  wire  _T_903 = _T_791 & REG_58; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_59; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_905 = 16'h1 << REG_59; // @[OneHot.scala 57:35]
  wire  _T_906 = waitInflightMask_13 == _T_905; // @[Sbuffer.scala 744:29]
  wire  _T_907 = _T_903 & _T_906; // @[Sbuffer.scala 743:30]
  reg  REG_60; // @[Sbuffer.scala 743:16]
  wire  _T_909 = _T_797 & REG_60; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_61; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_911 = 16'h1 << REG_61; // @[OneHot.scala 57:35]
  wire  _T_912 = waitInflightMask_14 == _T_911; // @[Sbuffer.scala 744:29]
  wire  _T_913 = _T_909 & _T_912; // @[Sbuffer.scala 743:30]
  reg  REG_62; // @[Sbuffer.scala 743:16]
  wire  _T_915 = _T_803 & REG_62; // @[Sbuffer.scala 742:33]
  reg [3:0] REG_63; // @[Sbuffer.scala 744:49]
  wire [15:0] _T_917 = 16'h1 << REG_63; // @[OneHot.scala 57:35]
  wire  _T_918 = waitInflightMask_15 == _T_917; // @[Sbuffer.scala 744:29]
  wire  _T_919 = _T_915 & _T_918; // @[Sbuffer.scala 743:30]
  wire [63:0] _dataModule_io_maskFlushReq_0_bits_wvec_T = 64'h1 << io_dcache_main_pipe_hit_resp_bits_id; // @[OneHot.scala 57:35]
  wire [63:0] _dataModule_io_maskFlushReq_1_bits_wvec_T = 64'h1 << io_dcache_refill_hit_resp_bits_id; // @[OneHot.scala 57:35]
  wire  _GEN_3164 = 4'h0 == io_dcache_replay_resp_bits_id[3:0] | _GEN_841; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3165 = 4'h1 == io_dcache_replay_resp_bits_id[3:0] | _GEN_842; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3166 = 4'h2 == io_dcache_replay_resp_bits_id[3:0] | _GEN_843; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3167 = 4'h3 == io_dcache_replay_resp_bits_id[3:0] | _GEN_844; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3168 = 4'h4 == io_dcache_replay_resp_bits_id[3:0] | _GEN_845; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3169 = 4'h5 == io_dcache_replay_resp_bits_id[3:0] | _GEN_846; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3170 = 4'h6 == io_dcache_replay_resp_bits_id[3:0] | _GEN_847; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3171 = 4'h7 == io_dcache_replay_resp_bits_id[3:0] | _GEN_848; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3172 = 4'h8 == io_dcache_replay_resp_bits_id[3:0] | _GEN_849; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3173 = 4'h9 == io_dcache_replay_resp_bits_id[3:0] | _GEN_850; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3174 = 4'ha == io_dcache_replay_resp_bits_id[3:0] | _GEN_851; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3175 = 4'hb == io_dcache_replay_resp_bits_id[3:0] | _GEN_852; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3176 = 4'hc == io_dcache_replay_resp_bits_id[3:0] | _GEN_853; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3177 = 4'hd == io_dcache_replay_resp_bits_id[3:0] | _GEN_854; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3178 = 4'he == io_dcache_replay_resp_bits_id[3:0] | _GEN_855; // @[Sbuffer.scala 760:{40,40}]
  wire  _GEN_3179 = 4'hf == io_dcache_replay_resp_bits_id[3:0] | _GEN_856; // @[Sbuffer.scala 760:{40,40}]
  wire [4:0] _missqReplayCount_0_T_1 = missqReplayCount_0 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_0_T_1 = cohCount_0 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_1_T_1 = missqReplayCount_1 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_1_T_1 = cohCount_1 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_2_T_1 = missqReplayCount_2 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_2_T_1 = cohCount_2 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_3_T_1 = missqReplayCount_3 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_3_T_1 = cohCount_3 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_4_T_1 = missqReplayCount_4 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_4_T_1 = cohCount_4 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_5_T_1 = missqReplayCount_5 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_5_T_1 = cohCount_5 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_6_T_1 = missqReplayCount_6 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_6_T_1 = cohCount_6 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_7_T_1 = missqReplayCount_7 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_7_T_1 = cohCount_7 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_8_T_1 = missqReplayCount_8 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_8_T_1 = cohCount_8 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_9_T_1 = missqReplayCount_9 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_9_T_1 = cohCount_9 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_10_T_1 = missqReplayCount_10 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_10_T_1 = cohCount_10 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_11_T_1 = missqReplayCount_11 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_11_T_1 = cohCount_11 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_12_T_1 = missqReplayCount_12 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_12_T_1 = cohCount_12 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_13_T_1 = missqReplayCount_13 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_13_T_1 = cohCount_13 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_14_T_1 = missqReplayCount_14 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_14_T_1 = cohCount_14 + 21'h1; // @[Sbuffer.scala 772:33]
  wire [4:0] _missqReplayCount_15_T_1 = missqReplayCount_15 + 5'h1; // @[Sbuffer.scala 769:50]
  wire [20:0] _cohCount_15_T_1 = cohCount_15 + 21'h1; // @[Sbuffer.scala 772:33]
  reg  tag_mismatch_REG; // @[Sbuffer.scala 799:31]
  reg  tag_mismatch_REG_31; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_30; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_31; // @[Reg.scala 19:16]
  wire  ptag_matches__15 = ptag_matches_r_30 == ptag_matches_r_31; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_32; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_47 = tag_mismatch_REG_31 != ptag_matches__15 & tag_mismatch_REG_32; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_29; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_28; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_29; // @[Reg.scala 19:16]
  wire  ptag_matches__14 = ptag_matches_r_28 == ptag_matches_r_29; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_30; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_44 = tag_mismatch_REG_29 != ptag_matches__14 & tag_mismatch_REG_30; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_27; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_26; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_27; // @[Reg.scala 19:16]
  wire  ptag_matches__13 = ptag_matches_r_26 == ptag_matches_r_27; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_28; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_41 = tag_mismatch_REG_27 != ptag_matches__13 & tag_mismatch_REG_28; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_25; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_24; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_25; // @[Reg.scala 19:16]
  wire  ptag_matches__12 = ptag_matches_r_24 == ptag_matches_r_25; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_26; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_38 = tag_mismatch_REG_25 != ptag_matches__12 & tag_mismatch_REG_26; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_23; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_22; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_23; // @[Reg.scala 19:16]
  wire  ptag_matches__11 = ptag_matches_r_22 == ptag_matches_r_23; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_24; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_35 = tag_mismatch_REG_23 != ptag_matches__11 & tag_mismatch_REG_24; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_21; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_20; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_21; // @[Reg.scala 19:16]
  wire  ptag_matches__10 = ptag_matches_r_20 == ptag_matches_r_21; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_22; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_32 = tag_mismatch_REG_21 != ptag_matches__10 & tag_mismatch_REG_22; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_19; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_18; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_19; // @[Reg.scala 19:16]
  wire  ptag_matches__9 = ptag_matches_r_18 == ptag_matches_r_19; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_20; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_29 = tag_mismatch_REG_19 != ptag_matches__9 & tag_mismatch_REG_20; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_17; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_16; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_17; // @[Reg.scala 19:16]
  wire  ptag_matches__8 = ptag_matches_r_16 == ptag_matches_r_17; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_18; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_26 = tag_mismatch_REG_17 != ptag_matches__8 & tag_mismatch_REG_18; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_15; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_14; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_15; // @[Reg.scala 19:16]
  wire  ptag_matches__7 = ptag_matches_r_14 == ptag_matches_r_15; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_16; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_23 = tag_mismatch_REG_15 != ptag_matches__7 & tag_mismatch_REG_16; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_13; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_12; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_13; // @[Reg.scala 19:16]
  wire  ptag_matches__6 = ptag_matches_r_12 == ptag_matches_r_13; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_14; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_20 = tag_mismatch_REG_13 != ptag_matches__6 & tag_mismatch_REG_14; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_11; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_10; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_11; // @[Reg.scala 19:16]
  wire  ptag_matches__5 = ptag_matches_r_10 == ptag_matches_r_11; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_12; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_17 = tag_mismatch_REG_11 != ptag_matches__5 & tag_mismatch_REG_12; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_9; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_8; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_9; // @[Reg.scala 19:16]
  wire  ptag_matches__4 = ptag_matches_r_8 == ptag_matches_r_9; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_10; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_14 = tag_mismatch_REG_9 != ptag_matches__4 & tag_mismatch_REG_10; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_7; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_6; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_7; // @[Reg.scala 19:16]
  wire  ptag_matches__3 = ptag_matches_r_6 == ptag_matches_r_7; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_8; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_11 = tag_mismatch_REG_7 != ptag_matches__3 & tag_mismatch_REG_8; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_5; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_4; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_5; // @[Reg.scala 19:16]
  wire  ptag_matches__2 = ptag_matches_r_4 == ptag_matches_r_5; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_6; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_8 = tag_mismatch_REG_5 != ptag_matches__2 & tag_mismatch_REG_6; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_3; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_2; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_3; // @[Reg.scala 19:16]
  wire  ptag_matches__1 = ptag_matches_r_2 == ptag_matches_r_3; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_4; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_5 = tag_mismatch_REG_3 != ptag_matches__1 & tag_mismatch_REG_4; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_1; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_1; // @[Reg.scala 19:16]
  wire  ptag_matches__0 = ptag_matches_r == ptag_matches_r_1; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_2; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_2 = tag_mismatch_REG_1 != ptag_matches__0 & tag_mismatch_REG_2; // @[Sbuffer.scala 800:52]
  wire [7:0] tag_mismatch_lo = {_tag_mismatch_T_23,_tag_mismatch_T_20,_tag_mismatch_T_17,_tag_mismatch_T_14,
    _tag_mismatch_T_11,_tag_mismatch_T_8,_tag_mismatch_T_5,_tag_mismatch_T_2}; // @[Sbuffer.scala 801:8]
  wire [15:0] _tag_mismatch_T_48 = {_tag_mismatch_T_47,_tag_mismatch_T_44,_tag_mismatch_T_41,_tag_mismatch_T_38,
    _tag_mismatch_T_35,_tag_mismatch_T_32,_tag_mismatch_T_29,_tag_mismatch_T_26,tag_mismatch_lo}; // @[Sbuffer.scala 801:8]
  wire  _tag_mismatch_T_49 = |_tag_mismatch_T_48; // @[Sbuffer.scala 801:15]
  wire  tag_mismatch = tag_mismatch_REG & _tag_mismatch_T_49; // @[Sbuffer.scala 799:47]
  reg  tag_mismatch_REG_33; // @[Sbuffer.scala 799:31]
  reg  tag_mismatch_REG_64; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_62; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_63; // @[Reg.scala 19:16]
  wire  ptag_matches_1_15 = ptag_matches_r_62 == ptag_matches_r_63; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_65; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_97 = tag_mismatch_REG_64 != ptag_matches_1_15 & tag_mismatch_REG_65; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_62; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_60; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_61; // @[Reg.scala 19:16]
  wire  ptag_matches_1_14 = ptag_matches_r_60 == ptag_matches_r_61; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_63; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_94 = tag_mismatch_REG_62 != ptag_matches_1_14 & tag_mismatch_REG_63; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_60; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_58; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_59; // @[Reg.scala 19:16]
  wire  ptag_matches_1_13 = ptag_matches_r_58 == ptag_matches_r_59; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_61; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_91 = tag_mismatch_REG_60 != ptag_matches_1_13 & tag_mismatch_REG_61; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_58; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_56; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_57; // @[Reg.scala 19:16]
  wire  ptag_matches_1_12 = ptag_matches_r_56 == ptag_matches_r_57; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_59; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_88 = tag_mismatch_REG_58 != ptag_matches_1_12 & tag_mismatch_REG_59; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_56; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_54; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_55; // @[Reg.scala 19:16]
  wire  ptag_matches_1_11 = ptag_matches_r_54 == ptag_matches_r_55; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_57; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_85 = tag_mismatch_REG_56 != ptag_matches_1_11 & tag_mismatch_REG_57; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_54; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_52; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_53; // @[Reg.scala 19:16]
  wire  ptag_matches_1_10 = ptag_matches_r_52 == ptag_matches_r_53; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_55; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_82 = tag_mismatch_REG_54 != ptag_matches_1_10 & tag_mismatch_REG_55; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_52; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_50; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_51; // @[Reg.scala 19:16]
  wire  ptag_matches_1_9 = ptag_matches_r_50 == ptag_matches_r_51; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_53; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_79 = tag_mismatch_REG_52 != ptag_matches_1_9 & tag_mismatch_REG_53; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_50; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_48; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_49; // @[Reg.scala 19:16]
  wire  ptag_matches_1_8 = ptag_matches_r_48 == ptag_matches_r_49; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_51; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_76 = tag_mismatch_REG_50 != ptag_matches_1_8 & tag_mismatch_REG_51; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_48; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_46; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_47; // @[Reg.scala 19:16]
  wire  ptag_matches_1_7 = ptag_matches_r_46 == ptag_matches_r_47; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_49; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_73 = tag_mismatch_REG_48 != ptag_matches_1_7 & tag_mismatch_REG_49; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_46; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_44; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_45; // @[Reg.scala 19:16]
  wire  ptag_matches_1_6 = ptag_matches_r_44 == ptag_matches_r_45; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_47; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_70 = tag_mismatch_REG_46 != ptag_matches_1_6 & tag_mismatch_REG_47; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_44; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_42; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_43; // @[Reg.scala 19:16]
  wire  ptag_matches_1_5 = ptag_matches_r_42 == ptag_matches_r_43; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_45; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_67 = tag_mismatch_REG_44 != ptag_matches_1_5 & tag_mismatch_REG_45; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_42; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_40; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_41; // @[Reg.scala 19:16]
  wire  ptag_matches_1_4 = ptag_matches_r_40 == ptag_matches_r_41; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_43; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_64 = tag_mismatch_REG_42 != ptag_matches_1_4 & tag_mismatch_REG_43; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_40; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_38; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_39; // @[Reg.scala 19:16]
  wire  ptag_matches_1_3 = ptag_matches_r_38 == ptag_matches_r_39; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_41; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_61 = tag_mismatch_REG_40 != ptag_matches_1_3 & tag_mismatch_REG_41; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_38; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_36; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_37; // @[Reg.scala 19:16]
  wire  ptag_matches_1_2 = ptag_matches_r_36 == ptag_matches_r_37; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_39; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_58 = tag_mismatch_REG_38 != ptag_matches_1_2 & tag_mismatch_REG_39; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_36; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_34; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_35; // @[Reg.scala 19:16]
  wire  ptag_matches_1_1 = ptag_matches_r_34 == ptag_matches_r_35; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_37; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_55 = tag_mismatch_REG_36 != ptag_matches_1_1 & tag_mismatch_REG_37; // @[Sbuffer.scala 800:52]
  reg  tag_mismatch_REG_34; // @[Sbuffer.scala 800:14]
  reg [29:0] ptag_matches_r_32; // @[Reg.scala 19:16]
  reg [29:0] ptag_matches_r_33; // @[Reg.scala 19:16]
  wire  ptag_matches_1_0 = ptag_matches_r_32 == ptag_matches_r_33; // @[Sbuffer.scala 797:80]
  reg  tag_mismatch_REG_35; // @[Sbuffer.scala 800:62]
  wire  _tag_mismatch_T_52 = tag_mismatch_REG_34 != ptag_matches_1_0 & tag_mismatch_REG_35; // @[Sbuffer.scala 800:52]
  wire [7:0] tag_mismatch_lo_1 = {_tag_mismatch_T_73,_tag_mismatch_T_70,_tag_mismatch_T_67,_tag_mismatch_T_64,
    _tag_mismatch_T_61,_tag_mismatch_T_58,_tag_mismatch_T_55,_tag_mismatch_T_52}; // @[Sbuffer.scala 801:8]
  wire [15:0] _tag_mismatch_T_98 = {_tag_mismatch_T_97,_tag_mismatch_T_94,_tag_mismatch_T_91,_tag_mismatch_T_88,
    _tag_mismatch_T_85,_tag_mismatch_T_82,_tag_mismatch_T_79,_tag_mismatch_T_76,tag_mismatch_lo_1}; // @[Sbuffer.scala 801:8]
  wire  _tag_mismatch_T_99 = |_tag_mismatch_T_98; // @[Sbuffer.scala 801:15]
  wire  tag_mismatch_1 = tag_mismatch_REG_33 & _tag_mismatch_T_99; // @[Sbuffer.scala 799:47]
  wire  vtag_matches__0 = vtag_0 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__1 = vtag_1 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__2 = vtag_2 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__3 = vtag_3 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__4 = vtag_4 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__5 = vtag_5 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__6 = vtag_6 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__7 = vtag_7 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__8 = vtag_8 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__9 = vtag_9 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__10 = vtag_10 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__11 = vtag_11 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__12 = vtag_12 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__13 = vtag_13 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__14 = vtag_14 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches__15 = vtag_15 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  reg  valid_tag_match_reg_0; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_2; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_3; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_4; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_5; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_6; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_7; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_8; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_9; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_10; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_11; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_12; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_13; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_14; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_15; // @[Sbuffer.scala 816:60]
  reg  inflight_tag_match_reg_0; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_2; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_3; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_4; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_5; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_6; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_7; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_8; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_9; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_10; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_11; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_12; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_13; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_14; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_15; // @[Sbuffer.scala 817:66]
  wire  _GEN_3294 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_0 : _GEN_1948; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3295 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_0 : _GEN_3294; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3296 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_0 : _GEN_3295; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3297 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_0 : _GEN_3296; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3302 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_1 : _GEN_1932; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3303 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_1 : _GEN_3302; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3304 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_1 : _GEN_3303; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3305 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_1 : _GEN_3304; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3310 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_2 : _GEN_1980; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3311 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_2 : _GEN_3310; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3312 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_2 : _GEN_3311; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3313 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_2 : _GEN_3312; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3318 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_3 : _GEN_1964; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3319 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_3 : _GEN_3318; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3320 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_3 : _GEN_3319; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3321 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_3 : _GEN_3320; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3326 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_4 : _GEN_2012; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3327 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_4 : _GEN_3326; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3328 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_4 : _GEN_3327; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3329 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_4 : _GEN_3328; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3334 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_5 : _GEN_1996; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3335 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_5 : _GEN_3334; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3336 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_5 : _GEN_3335; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3337 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_5 : _GEN_3336; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3342 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_6 : _GEN_2044; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3343 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_6 : _GEN_3342; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3344 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_6 : _GEN_3343; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3345 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_6 : _GEN_3344; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3350 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_1_7 : _GEN_2028; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3351 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_2_7 : _GEN_3350; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3352 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_3_7 : _GEN_3351; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3353 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_0_4_7 : _GEN_3352; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3358 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_0 : dataModule_io_maskOut_1_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3359 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_0 : _GEN_3358; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3360 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_0 : _GEN_3359; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3361 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_0 : _GEN_3360; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3366 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_1 : dataModule_io_maskOut_1_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3367 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_1 : _GEN_3366; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3368 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_1 : _GEN_3367; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3369 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_1 : _GEN_3368; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3374 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_2 : dataModule_io_maskOut_1_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3375 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_2 : _GEN_3374; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3376 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_2 : _GEN_3375; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3377 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_2 : _GEN_3376; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3382 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_3 : dataModule_io_maskOut_1_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3383 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_3 : _GEN_3382; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3384 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_3 : _GEN_3383; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3385 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_3 : _GEN_3384; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3390 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_4 : dataModule_io_maskOut_1_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3391 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_4 : _GEN_3390; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3392 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_4 : _GEN_3391; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3393 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_4 : _GEN_3392; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3398 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_5 : dataModule_io_maskOut_1_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3399 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_5 : _GEN_3398; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3400 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_5 : _GEN_3399; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3401 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_5 : _GEN_3400; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3406 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_6 : dataModule_io_maskOut_1_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3407 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_6 : _GEN_3406; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3408 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_6 : _GEN_3407; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3409 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_6 : _GEN_3408; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3414 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_1_7 : dataModule_io_maskOut_1_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3415 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_2_7 : _GEN_3414; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3416 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_3_7 : _GEN_3415; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3417 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_1_4_7 : _GEN_3416; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3422 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_0 : dataModule_io_maskOut_2_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3423 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_0 : _GEN_3422; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3424 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_0 : _GEN_3423; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3425 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_0 : _GEN_3424; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3430 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_1 : dataModule_io_maskOut_2_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3431 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_1 : _GEN_3430; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3432 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_1 : _GEN_3431; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3433 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_1 : _GEN_3432; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3438 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_2 : dataModule_io_maskOut_2_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3439 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_2 : _GEN_3438; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3440 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_2 : _GEN_3439; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3441 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_2 : _GEN_3440; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3446 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_3 : dataModule_io_maskOut_2_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3447 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_3 : _GEN_3446; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3448 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_3 : _GEN_3447; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3449 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_3 : _GEN_3448; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3454 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_4 : dataModule_io_maskOut_2_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3455 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_4 : _GEN_3454; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3456 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_4 : _GEN_3455; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3457 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_4 : _GEN_3456; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3462 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_5 : dataModule_io_maskOut_2_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3463 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_5 : _GEN_3462; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3464 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_5 : _GEN_3463; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3465 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_5 : _GEN_3464; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3470 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_6 : dataModule_io_maskOut_2_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3471 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_6 : _GEN_3470; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3472 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_6 : _GEN_3471; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3473 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_6 : _GEN_3472; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3478 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_1_7 : dataModule_io_maskOut_2_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3479 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_2_7 : _GEN_3478; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3480 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_3_7 : _GEN_3479; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3481 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_2_4_7 : _GEN_3480; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3486 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_0 : dataModule_io_maskOut_3_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3487 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_0 : _GEN_3486; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3488 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_0 : _GEN_3487; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3489 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_0 : _GEN_3488; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3494 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_1 : dataModule_io_maskOut_3_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3495 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_1 : _GEN_3494; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3496 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_1 : _GEN_3495; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3497 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_1 : _GEN_3496; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3502 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_2 : dataModule_io_maskOut_3_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3503 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_2 : _GEN_3502; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3504 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_2 : _GEN_3503; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3505 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_2 : _GEN_3504; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3510 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_3 : dataModule_io_maskOut_3_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3511 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_3 : _GEN_3510; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3512 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_3 : _GEN_3511; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3513 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_3 : _GEN_3512; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3518 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_4 : dataModule_io_maskOut_3_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3519 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_4 : _GEN_3518; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3520 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_4 : _GEN_3519; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3521 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_4 : _GEN_3520; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3526 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_5 : dataModule_io_maskOut_3_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3527 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_5 : _GEN_3526; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3528 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_5 : _GEN_3527; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3529 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_5 : _GEN_3528; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3534 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_6 : dataModule_io_maskOut_3_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3535 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_6 : _GEN_3534; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3536 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_6 : _GEN_3535; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3537 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_6 : _GEN_3536; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3542 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_1_7 : dataModule_io_maskOut_3_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3543 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_2_7 : _GEN_3542; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3544 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_3_7 : _GEN_3543; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3545 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_3_4_7 : _GEN_3544; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3550 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_0 : dataModule_io_maskOut_4_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3551 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_0 : _GEN_3550; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3552 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_0 : _GEN_3551; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3553 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_0 : _GEN_3552; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3558 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_1 : dataModule_io_maskOut_4_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3559 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_1 : _GEN_3558; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3560 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_1 : _GEN_3559; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3561 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_1 : _GEN_3560; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3566 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_2 : dataModule_io_maskOut_4_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3567 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_2 : _GEN_3566; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3568 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_2 : _GEN_3567; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3569 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_2 : _GEN_3568; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3574 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_3 : dataModule_io_maskOut_4_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3575 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_3 : _GEN_3574; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3576 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_3 : _GEN_3575; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3577 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_3 : _GEN_3576; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3582 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_4 : dataModule_io_maskOut_4_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3583 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_4 : _GEN_3582; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3584 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_4 : _GEN_3583; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3585 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_4 : _GEN_3584; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3590 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_5 : dataModule_io_maskOut_4_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3591 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_5 : _GEN_3590; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3592 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_5 : _GEN_3591; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3593 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_5 : _GEN_3592; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3598 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_6 : dataModule_io_maskOut_4_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3599 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_6 : _GEN_3598; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3600 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_6 : _GEN_3599; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3601 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_6 : _GEN_3600; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3606 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_1_7 : dataModule_io_maskOut_4_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3607 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_2_7 : _GEN_3606; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3608 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_3_7 : _GEN_3607; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3609 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_4_4_7 : _GEN_3608; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3614 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_0 : dataModule_io_maskOut_5_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3615 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_0 : _GEN_3614; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3616 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_0 : _GEN_3615; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3617 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_0 : _GEN_3616; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3622 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_1 : dataModule_io_maskOut_5_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3623 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_1 : _GEN_3622; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3624 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_1 : _GEN_3623; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3625 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_1 : _GEN_3624; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3630 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_2 : dataModule_io_maskOut_5_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3631 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_2 : _GEN_3630; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3632 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_2 : _GEN_3631; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3633 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_2 : _GEN_3632; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3638 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_3 : dataModule_io_maskOut_5_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3639 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_3 : _GEN_3638; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3640 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_3 : _GEN_3639; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3641 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_3 : _GEN_3640; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3646 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_4 : dataModule_io_maskOut_5_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3647 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_4 : _GEN_3646; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3648 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_4 : _GEN_3647; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3649 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_4 : _GEN_3648; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3654 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_5 : dataModule_io_maskOut_5_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3655 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_5 : _GEN_3654; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3656 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_5 : _GEN_3655; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3657 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_5 : _GEN_3656; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3662 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_6 : dataModule_io_maskOut_5_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3663 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_6 : _GEN_3662; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3664 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_6 : _GEN_3663; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3665 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_6 : _GEN_3664; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3670 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_1_7 : dataModule_io_maskOut_5_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3671 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_2_7 : _GEN_3670; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3672 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_3_7 : _GEN_3671; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3673 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_5_4_7 : _GEN_3672; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3678 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_0 : dataModule_io_maskOut_6_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3679 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_0 : _GEN_3678; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3680 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_0 : _GEN_3679; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3681 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_0 : _GEN_3680; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3686 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_1 : dataModule_io_maskOut_6_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3687 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_1 : _GEN_3686; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3688 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_1 : _GEN_3687; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3689 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_1 : _GEN_3688; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3694 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_2 : dataModule_io_maskOut_6_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3695 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_2 : _GEN_3694; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3696 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_2 : _GEN_3695; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3697 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_2 : _GEN_3696; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3702 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_3 : dataModule_io_maskOut_6_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3703 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_3 : _GEN_3702; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3704 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_3 : _GEN_3703; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3705 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_3 : _GEN_3704; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3710 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_4 : dataModule_io_maskOut_6_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3711 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_4 : _GEN_3710; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3712 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_4 : _GEN_3711; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3713 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_4 : _GEN_3712; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3718 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_5 : dataModule_io_maskOut_6_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3719 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_5 : _GEN_3718; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3720 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_5 : _GEN_3719; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3721 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_5 : _GEN_3720; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3726 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_6 : dataModule_io_maskOut_6_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3727 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_6 : _GEN_3726; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3728 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_6 : _GEN_3727; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3729 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_6 : _GEN_3728; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3734 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_1_7 : dataModule_io_maskOut_6_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3735 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_2_7 : _GEN_3734; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3736 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_3_7 : _GEN_3735; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3737 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_6_4_7 : _GEN_3736; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3742 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_0 : dataModule_io_maskOut_7_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3743 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_0 : _GEN_3742; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3744 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_0 : _GEN_3743; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3745 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_0 : _GEN_3744; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3750 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_1 : dataModule_io_maskOut_7_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3751 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_1 : _GEN_3750; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3752 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_1 : _GEN_3751; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3753 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_1 : _GEN_3752; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3758 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_2 : dataModule_io_maskOut_7_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3759 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_2 : _GEN_3758; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3760 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_2 : _GEN_3759; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3761 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_2 : _GEN_3760; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3766 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_3 : dataModule_io_maskOut_7_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3767 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_3 : _GEN_3766; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3768 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_3 : _GEN_3767; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3769 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_3 : _GEN_3768; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3774 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_4 : dataModule_io_maskOut_7_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3775 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_4 : _GEN_3774; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3776 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_4 : _GEN_3775; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3777 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_4 : _GEN_3776; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3782 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_5 : dataModule_io_maskOut_7_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3783 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_5 : _GEN_3782; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3784 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_5 : _GEN_3783; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3785 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_5 : _GEN_3784; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3790 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_6 : dataModule_io_maskOut_7_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3791 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_6 : _GEN_3790; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3792 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_6 : _GEN_3791; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3793 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_6 : _GEN_3792; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3798 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_1_7 : dataModule_io_maskOut_7_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3799 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_2_7 : _GEN_3798; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3800 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_3_7 : _GEN_3799; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3801 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_7_4_7 : _GEN_3800; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3806 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_0 : dataModule_io_maskOut_8_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3807 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_0 : _GEN_3806; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3808 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_0 : _GEN_3807; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3809 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_0 : _GEN_3808; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3814 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_1 : dataModule_io_maskOut_8_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3815 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_1 : _GEN_3814; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3816 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_1 : _GEN_3815; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3817 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_1 : _GEN_3816; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3822 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_2 : dataModule_io_maskOut_8_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3823 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_2 : _GEN_3822; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3824 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_2 : _GEN_3823; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3825 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_2 : _GEN_3824; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3830 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_3 : dataModule_io_maskOut_8_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3831 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_3 : _GEN_3830; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3832 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_3 : _GEN_3831; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3833 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_3 : _GEN_3832; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3838 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_4 : dataModule_io_maskOut_8_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3839 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_4 : _GEN_3838; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3840 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_4 : _GEN_3839; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3841 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_4 : _GEN_3840; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3846 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_5 : dataModule_io_maskOut_8_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3847 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_5 : _GEN_3846; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3848 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_5 : _GEN_3847; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3849 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_5 : _GEN_3848; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3854 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_6 : dataModule_io_maskOut_8_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3855 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_6 : _GEN_3854; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3856 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_6 : _GEN_3855; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3857 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_6 : _GEN_3856; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3862 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_1_7 : dataModule_io_maskOut_8_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3863 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_2_7 : _GEN_3862; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3864 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_3_7 : _GEN_3863; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3865 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_8_4_7 : _GEN_3864; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3870 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_0 : dataModule_io_maskOut_9_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3871 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_0 : _GEN_3870; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3872 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_0 : _GEN_3871; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3873 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_0 : _GEN_3872; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3878 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_1 : dataModule_io_maskOut_9_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3879 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_1 : _GEN_3878; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3880 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_1 : _GEN_3879; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3881 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_1 : _GEN_3880; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3886 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_2 : dataModule_io_maskOut_9_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3887 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_2 : _GEN_3886; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3888 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_2 : _GEN_3887; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3889 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_2 : _GEN_3888; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3894 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_3 : dataModule_io_maskOut_9_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3895 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_3 : _GEN_3894; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3896 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_3 : _GEN_3895; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3897 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_3 : _GEN_3896; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3902 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_4 : dataModule_io_maskOut_9_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3903 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_4 : _GEN_3902; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3904 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_4 : _GEN_3903; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3905 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_4 : _GEN_3904; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3910 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_5 : dataModule_io_maskOut_9_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3911 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_5 : _GEN_3910; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3912 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_5 : _GEN_3911; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3913 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_5 : _GEN_3912; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3918 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_6 : dataModule_io_maskOut_9_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3919 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_6 : _GEN_3918; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3920 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_6 : _GEN_3919; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3921 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_6 : _GEN_3920; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3926 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_1_7 : dataModule_io_maskOut_9_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3927 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_2_7 : _GEN_3926; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3928 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_3_7 : _GEN_3927; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3929 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_9_4_7 : _GEN_3928; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3934 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_0 : dataModule_io_maskOut_10_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3935 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_0 : _GEN_3934; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3936 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_0 : _GEN_3935; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3937 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_0 : _GEN_3936; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3942 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_1 : dataModule_io_maskOut_10_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3943 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_1 : _GEN_3942; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3944 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_1 : _GEN_3943; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3945 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_1 : _GEN_3944; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3950 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_2 : dataModule_io_maskOut_10_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3951 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_2 : _GEN_3950; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3952 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_2 : _GEN_3951; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3953 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_2 : _GEN_3952; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3958 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_3 : dataModule_io_maskOut_10_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3959 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_3 : _GEN_3958; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3960 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_3 : _GEN_3959; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3961 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_3 : _GEN_3960; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3966 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_4 : dataModule_io_maskOut_10_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3967 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_4 : _GEN_3966; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3968 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_4 : _GEN_3967; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3969 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_4 : _GEN_3968; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3974 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_5 : dataModule_io_maskOut_10_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3975 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_5 : _GEN_3974; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3976 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_5 : _GEN_3975; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3977 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_5 : _GEN_3976; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3982 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_6 : dataModule_io_maskOut_10_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3983 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_6 : _GEN_3982; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3984 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_6 : _GEN_3983; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3985 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_6 : _GEN_3984; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3990 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_1_7 : dataModule_io_maskOut_10_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3991 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_2_7 : _GEN_3990; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3992 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_3_7 : _GEN_3991; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3993 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_10_4_7 : _GEN_3992; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3998 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_0 : dataModule_io_maskOut_11_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_3999 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_0 : _GEN_3998; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4000 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_0 : _GEN_3999; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4001 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_0 : _GEN_4000; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4006 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_1 : dataModule_io_maskOut_11_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4007 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_1 : _GEN_4006; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4008 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_1 : _GEN_4007; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4009 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_1 : _GEN_4008; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4014 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_2 : dataModule_io_maskOut_11_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4015 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_2 : _GEN_4014; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4016 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_2 : _GEN_4015; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4017 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_2 : _GEN_4016; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4022 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_3 : dataModule_io_maskOut_11_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4023 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_3 : _GEN_4022; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4024 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_3 : _GEN_4023; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4025 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_3 : _GEN_4024; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4030 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_4 : dataModule_io_maskOut_11_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4031 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_4 : _GEN_4030; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4032 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_4 : _GEN_4031; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4033 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_4 : _GEN_4032; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4038 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_5 : dataModule_io_maskOut_11_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4039 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_5 : _GEN_4038; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4040 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_5 : _GEN_4039; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4041 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_5 : _GEN_4040; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4046 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_6 : dataModule_io_maskOut_11_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4047 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_6 : _GEN_4046; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4048 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_6 : _GEN_4047; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4049 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_6 : _GEN_4048; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4054 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_1_7 : dataModule_io_maskOut_11_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4055 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_2_7 : _GEN_4054; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4056 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_3_7 : _GEN_4055; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4057 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_11_4_7 : _GEN_4056; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4062 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_0 : dataModule_io_maskOut_12_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4063 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_0 : _GEN_4062; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4064 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_0 : _GEN_4063; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4065 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_0 : _GEN_4064; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4070 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_1 : dataModule_io_maskOut_12_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4071 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_1 : _GEN_4070; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4072 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_1 : _GEN_4071; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4073 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_1 : _GEN_4072; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4078 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_2 : dataModule_io_maskOut_12_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4079 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_2 : _GEN_4078; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4080 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_2 : _GEN_4079; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4081 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_2 : _GEN_4080; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4086 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_3 : dataModule_io_maskOut_12_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4087 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_3 : _GEN_4086; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4088 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_3 : _GEN_4087; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4089 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_3 : _GEN_4088; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4094 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_4 : dataModule_io_maskOut_12_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4095 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_4 : _GEN_4094; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4096 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_4 : _GEN_4095; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4097 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_4 : _GEN_4096; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4102 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_5 : dataModule_io_maskOut_12_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4103 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_5 : _GEN_4102; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4104 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_5 : _GEN_4103; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4105 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_5 : _GEN_4104; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4110 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_6 : dataModule_io_maskOut_12_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4111 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_6 : _GEN_4110; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4112 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_6 : _GEN_4111; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4113 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_6 : _GEN_4112; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4118 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_1_7 : dataModule_io_maskOut_12_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4119 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_2_7 : _GEN_4118; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4120 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_3_7 : _GEN_4119; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4121 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_12_4_7 : _GEN_4120; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4126 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_0 : dataModule_io_maskOut_13_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4127 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_0 : _GEN_4126; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4128 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_0 : _GEN_4127; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4129 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_0 : _GEN_4128; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4134 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_1 : dataModule_io_maskOut_13_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4135 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_1 : _GEN_4134; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4136 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_1 : _GEN_4135; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4137 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_1 : _GEN_4136; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4142 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_2 : dataModule_io_maskOut_13_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4143 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_2 : _GEN_4142; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4144 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_2 : _GEN_4143; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4145 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_2 : _GEN_4144; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4150 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_3 : dataModule_io_maskOut_13_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4151 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_3 : _GEN_4150; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4152 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_3 : _GEN_4151; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4153 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_3 : _GEN_4152; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4158 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_4 : dataModule_io_maskOut_13_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4159 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_4 : _GEN_4158; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4160 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_4 : _GEN_4159; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4161 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_4 : _GEN_4160; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4166 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_5 : dataModule_io_maskOut_13_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4167 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_5 : _GEN_4166; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4168 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_5 : _GEN_4167; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4169 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_5 : _GEN_4168; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4174 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_6 : dataModule_io_maskOut_13_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4175 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_6 : _GEN_4174; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4176 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_6 : _GEN_4175; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4177 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_6 : _GEN_4176; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4182 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_1_7 : dataModule_io_maskOut_13_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4183 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_2_7 : _GEN_4182; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4184 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_3_7 : _GEN_4183; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4185 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_13_4_7 : _GEN_4184; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4190 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_0 : dataModule_io_maskOut_14_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4191 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_0 : _GEN_4190; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4192 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_0 : _GEN_4191; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4193 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_0 : _GEN_4192; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4198 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_1 : dataModule_io_maskOut_14_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4199 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_1 : _GEN_4198; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4200 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_1 : _GEN_4199; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4201 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_1 : _GEN_4200; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4206 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_2 : dataModule_io_maskOut_14_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4207 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_2 : _GEN_4206; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4208 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_2 : _GEN_4207; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4209 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_2 : _GEN_4208; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4214 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_3 : dataModule_io_maskOut_14_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4215 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_3 : _GEN_4214; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4216 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_3 : _GEN_4215; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4217 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_3 : _GEN_4216; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4222 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_4 : dataModule_io_maskOut_14_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4223 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_4 : _GEN_4222; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4224 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_4 : _GEN_4223; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4225 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_4 : _GEN_4224; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4230 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_5 : dataModule_io_maskOut_14_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4231 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_5 : _GEN_4230; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4232 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_5 : _GEN_4231; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4233 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_5 : _GEN_4232; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4238 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_6 : dataModule_io_maskOut_14_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4239 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_6 : _GEN_4238; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4240 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_6 : _GEN_4239; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4241 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_6 : _GEN_4240; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4246 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_1_7 : dataModule_io_maskOut_14_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4247 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_2_7 : _GEN_4246; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4248 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_3_7 : _GEN_4247; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4249 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_14_4_7 : _GEN_4248; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4254 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_0 : dataModule_io_maskOut_15_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4255 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_0 : _GEN_4254; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4256 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_0 : _GEN_4255; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4257 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_0 : _GEN_4256; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4262 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_1 : dataModule_io_maskOut_15_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4263 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_1 : _GEN_4262; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4264 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_1 : _GEN_4263; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4265 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_1 : _GEN_4264; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4270 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_2 : dataModule_io_maskOut_15_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4271 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_2 : _GEN_4270; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4272 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_2 : _GEN_4271; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4273 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_2 : _GEN_4272; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4278 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_3 : dataModule_io_maskOut_15_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4279 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_3 : _GEN_4278; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4280 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_3 : _GEN_4279; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4281 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_3 : _GEN_4280; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4286 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_4 : dataModule_io_maskOut_15_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4287 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_4 : _GEN_4286; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4288 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_4 : _GEN_4287; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4289 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_4 : _GEN_4288; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4294 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_5 : dataModule_io_maskOut_15_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4295 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_5 : _GEN_4294; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4296 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_5 : _GEN_4295; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4297 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_5 : _GEN_4296; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4302 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_6 : dataModule_io_maskOut_15_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4303 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_6 : _GEN_4302; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4304 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_6 : _GEN_4303; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4305 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_6 : _GEN_4304; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4310 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_1_7 : dataModule_io_maskOut_15_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4311 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_2_7 : _GEN_4310; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4312 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_3_7 : _GEN_4311; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_4313 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_maskOut_15_4_7 : _GEN_4312; // @[Sbuffer.scala 820:{14,14}]
  reg  forward_mask_candidate_reg__0_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__0_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__1_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__2_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__3_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__4_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__5_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__6_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__7_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__8_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__9_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__10_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__11_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__12_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__13_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__14_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg__15_7; // @[Reg.scala 19:16]
  wire [7:0] _GEN_4446 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_0 : _GEN_924; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4447 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_0 : _GEN_4446; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4448 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_0 : _GEN_4447; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4449 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_0 : _GEN_4448; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4454 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_1 : _GEN_908; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4455 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_1 : _GEN_4454; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4456 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_1 : _GEN_4455; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4457 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_1 : _GEN_4456; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4462 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_2 : _GEN_956; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4463 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_2 : _GEN_4462; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4464 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_2 : _GEN_4463; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4465 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_2 : _GEN_4464; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4470 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_3 : _GEN_940; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4471 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_3 : _GEN_4470; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4472 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_3 : _GEN_4471; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4473 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_3 : _GEN_4472; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4478 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_4 : _GEN_988; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4479 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_4 : _GEN_4478; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4480 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_4 : _GEN_4479; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4481 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_4 : _GEN_4480; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4486 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_5 : _GEN_972; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4487 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_5 : _GEN_4486; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4488 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_5 : _GEN_4487; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4489 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_5 : _GEN_4488; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4494 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_6 : _GEN_1020; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4495 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_6 : _GEN_4494; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4496 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_6 : _GEN_4495; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4497 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_6 : _GEN_4496; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4502 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_1_7 : _GEN_1004; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4503 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_2_7 : _GEN_4502; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4504 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_3_7 : _GEN_4503; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4505 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_0_4_7 : _GEN_4504; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4509 = dataModule_io_dataOut_1_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4510 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_0 : _GEN_4509; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4511 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_0 : _GEN_4510; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4512 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_0 : _GEN_4511; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4513 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_0 : _GEN_4512; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4517 = dataModule_io_dataOut_1_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4518 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_1 : _GEN_4517; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4519 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_1 : _GEN_4518; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4520 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_1 : _GEN_4519; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4521 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_1 : _GEN_4520; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4525 = dataModule_io_dataOut_1_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4526 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_2 : _GEN_4525; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4527 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_2 : _GEN_4526; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4528 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_2 : _GEN_4527; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4529 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_2 : _GEN_4528; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4533 = dataModule_io_dataOut_1_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4534 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_3 : _GEN_4533; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4535 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_3 : _GEN_4534; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4536 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_3 : _GEN_4535; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4537 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_3 : _GEN_4536; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4541 = dataModule_io_dataOut_1_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4542 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_4 : _GEN_4541; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4543 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_4 : _GEN_4542; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4544 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_4 : _GEN_4543; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4545 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_4 : _GEN_4544; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4549 = dataModule_io_dataOut_1_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4550 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_5 : _GEN_4549; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4551 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_5 : _GEN_4550; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4552 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_5 : _GEN_4551; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4553 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_5 : _GEN_4552; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4557 = dataModule_io_dataOut_1_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4558 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_6 : _GEN_4557; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4559 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_6 : _GEN_4558; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4560 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_6 : _GEN_4559; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4561 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_6 : _GEN_4560; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4565 = dataModule_io_dataOut_1_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4566 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_1_7 : _GEN_4565; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4567 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_2_7 : _GEN_4566; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4568 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_3_7 : _GEN_4567; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4569 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_1_4_7 : _GEN_4568; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4573 = dataModule_io_dataOut_2_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4574 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_0 : _GEN_4573; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4575 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_0 : _GEN_4574; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4576 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_0 : _GEN_4575; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4577 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_0 : _GEN_4576; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4581 = dataModule_io_dataOut_2_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4582 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_1 : _GEN_4581; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4583 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_1 : _GEN_4582; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4584 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_1 : _GEN_4583; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4585 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_1 : _GEN_4584; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4589 = dataModule_io_dataOut_2_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4590 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_2 : _GEN_4589; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4591 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_2 : _GEN_4590; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4592 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_2 : _GEN_4591; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4593 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_2 : _GEN_4592; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4597 = dataModule_io_dataOut_2_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4598 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_3 : _GEN_4597; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4599 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_3 : _GEN_4598; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4600 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_3 : _GEN_4599; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4601 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_3 : _GEN_4600; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4605 = dataModule_io_dataOut_2_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4606 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_4 : _GEN_4605; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4607 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_4 : _GEN_4606; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4608 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_4 : _GEN_4607; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4609 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_4 : _GEN_4608; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4613 = dataModule_io_dataOut_2_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4614 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_5 : _GEN_4613; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4615 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_5 : _GEN_4614; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4616 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_5 : _GEN_4615; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4617 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_5 : _GEN_4616; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4621 = dataModule_io_dataOut_2_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4622 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_6 : _GEN_4621; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4623 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_6 : _GEN_4622; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4624 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_6 : _GEN_4623; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4625 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_6 : _GEN_4624; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4629 = dataModule_io_dataOut_2_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4630 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_1_7 : _GEN_4629; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4631 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_2_7 : _GEN_4630; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4632 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_3_7 : _GEN_4631; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4633 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_2_4_7 : _GEN_4632; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4637 = dataModule_io_dataOut_3_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4638 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_0 : _GEN_4637; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4639 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_0 : _GEN_4638; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4640 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_0 : _GEN_4639; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4641 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_0 : _GEN_4640; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4645 = dataModule_io_dataOut_3_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4646 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_1 : _GEN_4645; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4647 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_1 : _GEN_4646; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4648 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_1 : _GEN_4647; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4649 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_1 : _GEN_4648; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4653 = dataModule_io_dataOut_3_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4654 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_2 : _GEN_4653; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4655 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_2 : _GEN_4654; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4656 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_2 : _GEN_4655; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4657 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_2 : _GEN_4656; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4661 = dataModule_io_dataOut_3_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4662 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_3 : _GEN_4661; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4663 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_3 : _GEN_4662; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4664 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_3 : _GEN_4663; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4665 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_3 : _GEN_4664; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4669 = dataModule_io_dataOut_3_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4670 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_4 : _GEN_4669; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4671 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_4 : _GEN_4670; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4672 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_4 : _GEN_4671; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4673 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_4 : _GEN_4672; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4677 = dataModule_io_dataOut_3_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4678 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_5 : _GEN_4677; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4679 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_5 : _GEN_4678; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4680 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_5 : _GEN_4679; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4681 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_5 : _GEN_4680; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4685 = dataModule_io_dataOut_3_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4686 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_6 : _GEN_4685; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4687 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_6 : _GEN_4686; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4688 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_6 : _GEN_4687; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4689 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_6 : _GEN_4688; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4693 = dataModule_io_dataOut_3_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4694 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_1_7 : _GEN_4693; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4695 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_2_7 : _GEN_4694; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4696 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_3_7 : _GEN_4695; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4697 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_3_4_7 : _GEN_4696; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4701 = dataModule_io_dataOut_4_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4702 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_0 : _GEN_4701; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4703 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_0 : _GEN_4702; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4704 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_0 : _GEN_4703; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4705 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_0 : _GEN_4704; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4709 = dataModule_io_dataOut_4_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4710 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_1 : _GEN_4709; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4711 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_1 : _GEN_4710; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4712 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_1 : _GEN_4711; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4713 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_1 : _GEN_4712; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4717 = dataModule_io_dataOut_4_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4718 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_2 : _GEN_4717; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4719 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_2 : _GEN_4718; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4720 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_2 : _GEN_4719; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4721 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_2 : _GEN_4720; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4725 = dataModule_io_dataOut_4_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4726 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_3 : _GEN_4725; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4727 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_3 : _GEN_4726; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4728 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_3 : _GEN_4727; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4729 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_3 : _GEN_4728; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4733 = dataModule_io_dataOut_4_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4734 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_4 : _GEN_4733; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4735 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_4 : _GEN_4734; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4736 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_4 : _GEN_4735; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4737 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_4 : _GEN_4736; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4741 = dataModule_io_dataOut_4_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4742 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_5 : _GEN_4741; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4743 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_5 : _GEN_4742; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4744 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_5 : _GEN_4743; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4745 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_5 : _GEN_4744; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4749 = dataModule_io_dataOut_4_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4750 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_6 : _GEN_4749; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4751 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_6 : _GEN_4750; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4752 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_6 : _GEN_4751; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4753 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_6 : _GEN_4752; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4757 = dataModule_io_dataOut_4_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4758 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_1_7 : _GEN_4757; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4759 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_2_7 : _GEN_4758; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4760 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_3_7 : _GEN_4759; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4761 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_4_4_7 : _GEN_4760; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4765 = dataModule_io_dataOut_5_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4766 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_0 : _GEN_4765; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4767 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_0 : _GEN_4766; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4768 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_0 : _GEN_4767; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4769 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_0 : _GEN_4768; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4773 = dataModule_io_dataOut_5_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4774 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_1 : _GEN_4773; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4775 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_1 : _GEN_4774; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4776 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_1 : _GEN_4775; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4777 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_1 : _GEN_4776; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4781 = dataModule_io_dataOut_5_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4782 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_2 : _GEN_4781; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4783 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_2 : _GEN_4782; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4784 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_2 : _GEN_4783; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4785 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_2 : _GEN_4784; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4789 = dataModule_io_dataOut_5_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4790 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_3 : _GEN_4789; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4791 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_3 : _GEN_4790; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4792 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_3 : _GEN_4791; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4793 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_3 : _GEN_4792; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4797 = dataModule_io_dataOut_5_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4798 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_4 : _GEN_4797; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4799 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_4 : _GEN_4798; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4800 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_4 : _GEN_4799; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4801 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_4 : _GEN_4800; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4805 = dataModule_io_dataOut_5_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4806 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_5 : _GEN_4805; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4807 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_5 : _GEN_4806; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4808 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_5 : _GEN_4807; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4809 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_5 : _GEN_4808; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4813 = dataModule_io_dataOut_5_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4814 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_6 : _GEN_4813; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4815 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_6 : _GEN_4814; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4816 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_6 : _GEN_4815; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4817 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_6 : _GEN_4816; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4821 = dataModule_io_dataOut_5_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4822 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_1_7 : _GEN_4821; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4823 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_2_7 : _GEN_4822; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4824 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_3_7 : _GEN_4823; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4825 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_5_4_7 : _GEN_4824; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4829 = dataModule_io_dataOut_6_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4830 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_0 : _GEN_4829; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4831 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_0 : _GEN_4830; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4832 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_0 : _GEN_4831; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4833 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_0 : _GEN_4832; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4837 = dataModule_io_dataOut_6_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4838 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_1 : _GEN_4837; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4839 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_1 : _GEN_4838; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4840 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_1 : _GEN_4839; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4841 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_1 : _GEN_4840; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4845 = dataModule_io_dataOut_6_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4846 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_2 : _GEN_4845; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4847 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_2 : _GEN_4846; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4848 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_2 : _GEN_4847; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4849 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_2 : _GEN_4848; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4853 = dataModule_io_dataOut_6_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4854 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_3 : _GEN_4853; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4855 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_3 : _GEN_4854; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4856 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_3 : _GEN_4855; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4857 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_3 : _GEN_4856; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4861 = dataModule_io_dataOut_6_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4862 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_4 : _GEN_4861; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4863 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_4 : _GEN_4862; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4864 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_4 : _GEN_4863; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4865 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_4 : _GEN_4864; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4869 = dataModule_io_dataOut_6_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4870 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_5 : _GEN_4869; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4871 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_5 : _GEN_4870; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4872 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_5 : _GEN_4871; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4873 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_5 : _GEN_4872; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4877 = dataModule_io_dataOut_6_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4878 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_6 : _GEN_4877; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4879 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_6 : _GEN_4878; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4880 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_6 : _GEN_4879; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4881 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_6 : _GEN_4880; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4885 = dataModule_io_dataOut_6_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4886 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_1_7 : _GEN_4885; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4887 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_2_7 : _GEN_4886; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4888 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_3_7 : _GEN_4887; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4889 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_6_4_7 : _GEN_4888; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4893 = dataModule_io_dataOut_7_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4894 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_0 : _GEN_4893; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4895 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_0 : _GEN_4894; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4896 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_0 : _GEN_4895; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4897 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_0 : _GEN_4896; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4901 = dataModule_io_dataOut_7_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4902 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_1 : _GEN_4901; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4903 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_1 : _GEN_4902; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4904 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_1 : _GEN_4903; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4905 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_1 : _GEN_4904; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4909 = dataModule_io_dataOut_7_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4910 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_2 : _GEN_4909; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4911 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_2 : _GEN_4910; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4912 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_2 : _GEN_4911; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4913 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_2 : _GEN_4912; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4917 = dataModule_io_dataOut_7_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4918 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_3 : _GEN_4917; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4919 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_3 : _GEN_4918; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4920 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_3 : _GEN_4919; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4921 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_3 : _GEN_4920; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4925 = dataModule_io_dataOut_7_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4926 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_4 : _GEN_4925; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4927 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_4 : _GEN_4926; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4928 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_4 : _GEN_4927; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4929 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_4 : _GEN_4928; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4933 = dataModule_io_dataOut_7_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4934 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_5 : _GEN_4933; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4935 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_5 : _GEN_4934; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4936 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_5 : _GEN_4935; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4937 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_5 : _GEN_4936; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4941 = dataModule_io_dataOut_7_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4942 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_6 : _GEN_4941; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4943 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_6 : _GEN_4942; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4944 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_6 : _GEN_4943; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4945 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_6 : _GEN_4944; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4949 = dataModule_io_dataOut_7_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4950 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_1_7 : _GEN_4949; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4951 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_2_7 : _GEN_4950; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4952 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_3_7 : _GEN_4951; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4953 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_7_4_7 : _GEN_4952; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4957 = dataModule_io_dataOut_8_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4958 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_0 : _GEN_4957; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4959 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_0 : _GEN_4958; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4960 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_0 : _GEN_4959; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4961 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_0 : _GEN_4960; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4965 = dataModule_io_dataOut_8_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4966 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_1 : _GEN_4965; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4967 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_1 : _GEN_4966; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4968 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_1 : _GEN_4967; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4969 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_1 : _GEN_4968; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4973 = dataModule_io_dataOut_8_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4974 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_2 : _GEN_4973; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4975 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_2 : _GEN_4974; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4976 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_2 : _GEN_4975; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4977 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_2 : _GEN_4976; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4981 = dataModule_io_dataOut_8_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4982 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_3 : _GEN_4981; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4983 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_3 : _GEN_4982; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4984 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_3 : _GEN_4983; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4985 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_3 : _GEN_4984; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4989 = dataModule_io_dataOut_8_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4990 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_4 : _GEN_4989; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4991 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_4 : _GEN_4990; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4992 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_4 : _GEN_4991; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4993 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_4 : _GEN_4992; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4997 = dataModule_io_dataOut_8_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4998 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_5 : _GEN_4997; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_4999 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_5 : _GEN_4998; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5000 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_5 : _GEN_4999; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5001 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_5 : _GEN_5000; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5005 = dataModule_io_dataOut_8_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5006 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_6 : _GEN_5005; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5007 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_6 : _GEN_5006; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5008 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_6 : _GEN_5007; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5009 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_6 : _GEN_5008; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5013 = dataModule_io_dataOut_8_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5014 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_1_7 : _GEN_5013; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5015 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_2_7 : _GEN_5014; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5016 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_3_7 : _GEN_5015; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5017 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_8_4_7 : _GEN_5016; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5021 = dataModule_io_dataOut_9_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5022 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_0 : _GEN_5021; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5023 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_0 : _GEN_5022; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5024 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_0 : _GEN_5023; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5025 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_0 : _GEN_5024; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5029 = dataModule_io_dataOut_9_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5030 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_1 : _GEN_5029; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5031 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_1 : _GEN_5030; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5032 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_1 : _GEN_5031; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5033 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_1 : _GEN_5032; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5037 = dataModule_io_dataOut_9_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5038 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_2 : _GEN_5037; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5039 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_2 : _GEN_5038; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5040 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_2 : _GEN_5039; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5041 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_2 : _GEN_5040; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5045 = dataModule_io_dataOut_9_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5046 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_3 : _GEN_5045; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5047 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_3 : _GEN_5046; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5048 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_3 : _GEN_5047; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5049 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_3 : _GEN_5048; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5053 = dataModule_io_dataOut_9_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5054 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_4 : _GEN_5053; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5055 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_4 : _GEN_5054; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5056 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_4 : _GEN_5055; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5057 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_4 : _GEN_5056; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5061 = dataModule_io_dataOut_9_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5062 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_5 : _GEN_5061; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5063 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_5 : _GEN_5062; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5064 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_5 : _GEN_5063; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5065 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_5 : _GEN_5064; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5069 = dataModule_io_dataOut_9_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5070 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_6 : _GEN_5069; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5071 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_6 : _GEN_5070; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5072 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_6 : _GEN_5071; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5073 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_6 : _GEN_5072; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5077 = dataModule_io_dataOut_9_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5078 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_1_7 : _GEN_5077; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5079 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_2_7 : _GEN_5078; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5080 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_3_7 : _GEN_5079; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5081 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_9_4_7 : _GEN_5080; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5085 = dataModule_io_dataOut_10_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5086 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_0 : _GEN_5085; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5087 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_0 : _GEN_5086; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5088 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_0 : _GEN_5087; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5089 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_0 : _GEN_5088; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5093 = dataModule_io_dataOut_10_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5094 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_1 : _GEN_5093; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5095 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_1 : _GEN_5094; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5096 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_1 : _GEN_5095; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5097 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_1 : _GEN_5096; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5101 = dataModule_io_dataOut_10_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5102 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_2 : _GEN_5101; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5103 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_2 : _GEN_5102; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5104 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_2 : _GEN_5103; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5105 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_2 : _GEN_5104; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5109 = dataModule_io_dataOut_10_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5110 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_3 : _GEN_5109; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5111 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_3 : _GEN_5110; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5112 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_3 : _GEN_5111; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5113 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_3 : _GEN_5112; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5117 = dataModule_io_dataOut_10_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5118 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_4 : _GEN_5117; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5119 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_4 : _GEN_5118; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5120 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_4 : _GEN_5119; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5121 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_4 : _GEN_5120; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5125 = dataModule_io_dataOut_10_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5126 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_5 : _GEN_5125; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5127 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_5 : _GEN_5126; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5128 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_5 : _GEN_5127; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5129 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_5 : _GEN_5128; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5133 = dataModule_io_dataOut_10_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5134 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_6 : _GEN_5133; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5135 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_6 : _GEN_5134; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5136 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_6 : _GEN_5135; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5137 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_6 : _GEN_5136; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5141 = dataModule_io_dataOut_10_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5142 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_1_7 : _GEN_5141; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5143 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_2_7 : _GEN_5142; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5144 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_3_7 : _GEN_5143; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5145 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_10_4_7 : _GEN_5144; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5149 = dataModule_io_dataOut_11_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5150 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_0 : _GEN_5149; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5151 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_0 : _GEN_5150; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5152 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_0 : _GEN_5151; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5153 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_0 : _GEN_5152; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5157 = dataModule_io_dataOut_11_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5158 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_1 : _GEN_5157; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5159 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_1 : _GEN_5158; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5160 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_1 : _GEN_5159; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5161 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_1 : _GEN_5160; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5165 = dataModule_io_dataOut_11_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5166 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_2 : _GEN_5165; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5167 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_2 : _GEN_5166; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5168 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_2 : _GEN_5167; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5169 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_2 : _GEN_5168; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5173 = dataModule_io_dataOut_11_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5174 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_3 : _GEN_5173; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5175 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_3 : _GEN_5174; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5176 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_3 : _GEN_5175; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5177 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_3 : _GEN_5176; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5181 = dataModule_io_dataOut_11_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5182 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_4 : _GEN_5181; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5183 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_4 : _GEN_5182; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5184 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_4 : _GEN_5183; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5185 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_4 : _GEN_5184; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5189 = dataModule_io_dataOut_11_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5190 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_5 : _GEN_5189; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5191 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_5 : _GEN_5190; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5192 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_5 : _GEN_5191; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5193 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_5 : _GEN_5192; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5197 = dataModule_io_dataOut_11_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5198 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_6 : _GEN_5197; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5199 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_6 : _GEN_5198; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5200 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_6 : _GEN_5199; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5201 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_6 : _GEN_5200; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5205 = dataModule_io_dataOut_11_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5206 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_1_7 : _GEN_5205; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5207 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_2_7 : _GEN_5206; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5208 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_3_7 : _GEN_5207; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5209 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_11_4_7 : _GEN_5208; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5213 = dataModule_io_dataOut_12_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5214 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_0 : _GEN_5213; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5215 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_0 : _GEN_5214; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5216 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_0 : _GEN_5215; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5217 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_0 : _GEN_5216; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5221 = dataModule_io_dataOut_12_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5222 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_1 : _GEN_5221; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5223 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_1 : _GEN_5222; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5224 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_1 : _GEN_5223; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5225 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_1 : _GEN_5224; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5229 = dataModule_io_dataOut_12_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5230 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_2 : _GEN_5229; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5231 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_2 : _GEN_5230; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5232 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_2 : _GEN_5231; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5233 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_2 : _GEN_5232; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5237 = dataModule_io_dataOut_12_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5238 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_3 : _GEN_5237; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5239 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_3 : _GEN_5238; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5240 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_3 : _GEN_5239; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5241 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_3 : _GEN_5240; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5245 = dataModule_io_dataOut_12_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5246 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_4 : _GEN_5245; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5247 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_4 : _GEN_5246; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5248 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_4 : _GEN_5247; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5249 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_4 : _GEN_5248; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5253 = dataModule_io_dataOut_12_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5254 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_5 : _GEN_5253; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5255 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_5 : _GEN_5254; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5256 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_5 : _GEN_5255; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5257 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_5 : _GEN_5256; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5261 = dataModule_io_dataOut_12_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5262 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_6 : _GEN_5261; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5263 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_6 : _GEN_5262; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5264 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_6 : _GEN_5263; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5265 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_6 : _GEN_5264; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5269 = dataModule_io_dataOut_12_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5270 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_1_7 : _GEN_5269; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5271 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_2_7 : _GEN_5270; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5272 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_3_7 : _GEN_5271; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5273 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_12_4_7 : _GEN_5272; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5277 = dataModule_io_dataOut_13_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5278 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_0 : _GEN_5277; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5279 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_0 : _GEN_5278; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5280 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_0 : _GEN_5279; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5281 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_0 : _GEN_5280; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5285 = dataModule_io_dataOut_13_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5286 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_1 : _GEN_5285; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5287 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_1 : _GEN_5286; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5288 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_1 : _GEN_5287; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5289 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_1 : _GEN_5288; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5293 = dataModule_io_dataOut_13_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5294 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_2 : _GEN_5293; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5295 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_2 : _GEN_5294; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5296 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_2 : _GEN_5295; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5297 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_2 : _GEN_5296; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5301 = dataModule_io_dataOut_13_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5302 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_3 : _GEN_5301; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5303 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_3 : _GEN_5302; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5304 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_3 : _GEN_5303; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5305 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_3 : _GEN_5304; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5309 = dataModule_io_dataOut_13_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5310 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_4 : _GEN_5309; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5311 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_4 : _GEN_5310; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5312 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_4 : _GEN_5311; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5313 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_4 : _GEN_5312; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5317 = dataModule_io_dataOut_13_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5318 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_5 : _GEN_5317; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5319 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_5 : _GEN_5318; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5320 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_5 : _GEN_5319; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5321 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_5 : _GEN_5320; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5325 = dataModule_io_dataOut_13_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5326 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_6 : _GEN_5325; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5327 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_6 : _GEN_5326; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5328 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_6 : _GEN_5327; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5329 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_6 : _GEN_5328; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5333 = dataModule_io_dataOut_13_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5334 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_1_7 : _GEN_5333; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5335 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_2_7 : _GEN_5334; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5336 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_3_7 : _GEN_5335; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5337 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_13_4_7 : _GEN_5336; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5341 = dataModule_io_dataOut_14_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5342 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_0 : _GEN_5341; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5343 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_0 : _GEN_5342; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5344 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_0 : _GEN_5343; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5345 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_0 : _GEN_5344; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5349 = dataModule_io_dataOut_14_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5350 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_1 : _GEN_5349; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5351 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_1 : _GEN_5350; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5352 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_1 : _GEN_5351; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5353 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_1 : _GEN_5352; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5357 = dataModule_io_dataOut_14_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5358 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_2 : _GEN_5357; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5359 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_2 : _GEN_5358; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5360 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_2 : _GEN_5359; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5361 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_2 : _GEN_5360; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5365 = dataModule_io_dataOut_14_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5366 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_3 : _GEN_5365; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5367 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_3 : _GEN_5366; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5368 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_3 : _GEN_5367; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5369 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_3 : _GEN_5368; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5373 = dataModule_io_dataOut_14_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5374 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_4 : _GEN_5373; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5375 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_4 : _GEN_5374; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5376 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_4 : _GEN_5375; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5377 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_4 : _GEN_5376; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5381 = dataModule_io_dataOut_14_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5382 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_5 : _GEN_5381; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5383 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_5 : _GEN_5382; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5384 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_5 : _GEN_5383; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5385 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_5 : _GEN_5384; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5389 = dataModule_io_dataOut_14_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5390 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_6 : _GEN_5389; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5391 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_6 : _GEN_5390; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5392 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_6 : _GEN_5391; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5393 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_6 : _GEN_5392; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5397 = dataModule_io_dataOut_14_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5398 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_1_7 : _GEN_5397; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5399 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_2_7 : _GEN_5398; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5400 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_3_7 : _GEN_5399; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5401 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_14_4_7 : _GEN_5400; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5405 = dataModule_io_dataOut_15_0_0; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5406 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_0 : _GEN_5405; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5407 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_0 : _GEN_5406; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5408 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_0 : _GEN_5407; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5409 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_0 : _GEN_5408; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5413 = dataModule_io_dataOut_15_0_1; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5414 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_1 : _GEN_5413; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5415 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_1 : _GEN_5414; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5416 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_1 : _GEN_5415; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5417 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_1 : _GEN_5416; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5421 = dataModule_io_dataOut_15_0_2; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5422 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_2 : _GEN_5421; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5423 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_2 : _GEN_5422; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5424 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_2 : _GEN_5423; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5425 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_2 : _GEN_5424; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5429 = dataModule_io_dataOut_15_0_3; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5430 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_3 : _GEN_5429; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5431 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_3 : _GEN_5430; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5432 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_3 : _GEN_5431; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5433 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_3 : _GEN_5432; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5437 = dataModule_io_dataOut_15_0_4; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5438 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_4 : _GEN_5437; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5439 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_4 : _GEN_5438; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5440 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_4 : _GEN_5439; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5441 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_4 : _GEN_5440; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5445 = dataModule_io_dataOut_15_0_5; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5446 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_5 : _GEN_5445; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5447 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_5 : _GEN_5446; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5448 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_5 : _GEN_5447; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5449 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_5 : _GEN_5448; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5453 = dataModule_io_dataOut_15_0_6; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5454 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_6 : _GEN_5453; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5455 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_6 : _GEN_5454; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5456 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_6 : _GEN_5455; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5457 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_6 : _GEN_5456; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5461 = dataModule_io_dataOut_15_0_7; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5462 = 3'h1 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_1_7 : _GEN_5461; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5463 = 3'h2 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_2_7 : _GEN_5462; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5464 = 3'h3 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_3_7 : _GEN_5463; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_5465 = 3'h4 == io_forward_0_paddr[5:3] ? dataModule_io_dataOut_15_4_7 : _GEN_5464; // @[Sbuffer.scala 824:{14,14}]
  reg [7:0] forward_data_candidate_reg__0_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__0_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__1_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__2_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__3_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__4_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__5_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__6_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__7_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__8_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__9_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__10_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__11_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__12_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__13_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__14_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg__15_7; // @[Reg.scala 19:16]
  wire  _selectedValidMask_T_15 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_0; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_0 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_0 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_0 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_0 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_0 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_0 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_0 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_0 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_0 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_0 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_0 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_0 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_0 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_0 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_0 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_0 | _selectedValidMask_T_15; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_46 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_1; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_1 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_1 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_1 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_1 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_1 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_1 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_1 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_1 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_1 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_1 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_1 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_1 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_1 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_1 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_1 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_1 | _selectedValidMask_T_46; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_77 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_2; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_2 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_2 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_2 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_2 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_2 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_2 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_2 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_2 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_2 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_2 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_2 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_2 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_2 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_2 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_2 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_2 | _selectedValidMask_T_77; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_108 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_3; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_3 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_3 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_3 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_3 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_3 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_3 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_3 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_3 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_3 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_3 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_3 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_3 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_3 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_3 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_3 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_3 | _selectedValidMask_T_108; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_139 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_4; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_4 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_4 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_4 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_4 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_4 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_4 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_4 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_4 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_4 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_4 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_4 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_4 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_4 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_4 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_4 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_4 | _selectedValidMask_T_139; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_170 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_5; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_5 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_5 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_5 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_5 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_5 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_5 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_5 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_5 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_5 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_5 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_5 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_5 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_5 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_5 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_5 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_5 | _selectedValidMask_T_170; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_201 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_6; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_6 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_6 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_6 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_6 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_6 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_6 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_6 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_6 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_6 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_6 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_6 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_6 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_6 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_6 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_6 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_6 | _selectedValidMask_T_201; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_232 = valid_tag_match_reg_15 & forward_mask_candidate_reg__15_7; // @[Mux.scala 27:73]
  wire  selectedValidMask_0_7 = valid_tag_match_reg_0 & forward_mask_candidate_reg__0_7 | valid_tag_match_reg_1 &
    forward_mask_candidate_reg__1_7 | valid_tag_match_reg_2 & forward_mask_candidate_reg__2_7 | valid_tag_match_reg_3 &
    forward_mask_candidate_reg__3_7 | valid_tag_match_reg_4 & forward_mask_candidate_reg__4_7 | valid_tag_match_reg_5 &
    forward_mask_candidate_reg__5_7 | valid_tag_match_reg_6 & forward_mask_candidate_reg__6_7 | valid_tag_match_reg_7 &
    forward_mask_candidate_reg__7_7 | valid_tag_match_reg_8 & forward_mask_candidate_reg__8_7 | valid_tag_match_reg_9 &
    forward_mask_candidate_reg__9_7 | valid_tag_match_reg_10 & forward_mask_candidate_reg__10_7 | valid_tag_match_reg_11
     & forward_mask_candidate_reg__11_7 | valid_tag_match_reg_12 & forward_mask_candidate_reg__12_7 |
    valid_tag_match_reg_13 & forward_mask_candidate_reg__13_7 | valid_tag_match_reg_14 &
    forward_mask_candidate_reg__14_7 | _selectedValidMask_T_232; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_1 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_2 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_3 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_4 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_5 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_6 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_7 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_8 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_9 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_10 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_11 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_12 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_13 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_14 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_15 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_16 = _selectedValidData_T | _selectedValidData_T_1; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_17 = _selectedValidData_T_16 | _selectedValidData_T_2; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_18 = _selectedValidData_T_17 | _selectedValidData_T_3; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_19 = _selectedValidData_T_18 | _selectedValidData_T_4; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_20 = _selectedValidData_T_19 | _selectedValidData_T_5; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_21 = _selectedValidData_T_20 | _selectedValidData_T_6; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_22 = _selectedValidData_T_21 | _selectedValidData_T_7; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_23 = _selectedValidData_T_22 | _selectedValidData_T_8; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_24 = _selectedValidData_T_23 | _selectedValidData_T_9; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_25 = _selectedValidData_T_24 | _selectedValidData_T_10; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_26 = _selectedValidData_T_25 | _selectedValidData_T_11; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_27 = _selectedValidData_T_26 | _selectedValidData_T_12; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_28 = _selectedValidData_T_27 | _selectedValidData_T_13; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_29 = _selectedValidData_T_28 | _selectedValidData_T_14; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_0 = _selectedValidData_T_29 | _selectedValidData_T_15; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_31 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_32 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_33 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_34 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_35 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_36 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_37 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_38 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_39 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_40 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_41 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_42 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_43 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_44 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_45 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_46 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_47 = _selectedValidData_T_31 | _selectedValidData_T_32; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_48 = _selectedValidData_T_47 | _selectedValidData_T_33; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_49 = _selectedValidData_T_48 | _selectedValidData_T_34; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_50 = _selectedValidData_T_49 | _selectedValidData_T_35; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_51 = _selectedValidData_T_50 | _selectedValidData_T_36; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_52 = _selectedValidData_T_51 | _selectedValidData_T_37; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_53 = _selectedValidData_T_52 | _selectedValidData_T_38; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_54 = _selectedValidData_T_53 | _selectedValidData_T_39; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_55 = _selectedValidData_T_54 | _selectedValidData_T_40; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_56 = _selectedValidData_T_55 | _selectedValidData_T_41; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_57 = _selectedValidData_T_56 | _selectedValidData_T_42; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_58 = _selectedValidData_T_57 | _selectedValidData_T_43; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_59 = _selectedValidData_T_58 | _selectedValidData_T_44; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_60 = _selectedValidData_T_59 | _selectedValidData_T_45; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_1 = _selectedValidData_T_60 | _selectedValidData_T_46; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_62 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_63 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_64 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_65 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_66 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_67 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_68 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_69 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_70 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_71 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_72 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_73 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_74 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_75 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_76 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_77 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_78 = _selectedValidData_T_62 | _selectedValidData_T_63; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_79 = _selectedValidData_T_78 | _selectedValidData_T_64; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_80 = _selectedValidData_T_79 | _selectedValidData_T_65; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_81 = _selectedValidData_T_80 | _selectedValidData_T_66; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_82 = _selectedValidData_T_81 | _selectedValidData_T_67; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_83 = _selectedValidData_T_82 | _selectedValidData_T_68; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_84 = _selectedValidData_T_83 | _selectedValidData_T_69; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_85 = _selectedValidData_T_84 | _selectedValidData_T_70; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_86 = _selectedValidData_T_85 | _selectedValidData_T_71; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_87 = _selectedValidData_T_86 | _selectedValidData_T_72; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_88 = _selectedValidData_T_87 | _selectedValidData_T_73; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_89 = _selectedValidData_T_88 | _selectedValidData_T_74; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_90 = _selectedValidData_T_89 | _selectedValidData_T_75; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_91 = _selectedValidData_T_90 | _selectedValidData_T_76; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_2 = _selectedValidData_T_91 | _selectedValidData_T_77; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_93 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_94 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_95 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_96 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_97 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_98 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_99 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_100 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_101 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_102 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_103 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_104 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_105 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_106 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_107 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_108 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_109 = _selectedValidData_T_93 | _selectedValidData_T_94; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_110 = _selectedValidData_T_109 | _selectedValidData_T_95; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_111 = _selectedValidData_T_110 | _selectedValidData_T_96; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_112 = _selectedValidData_T_111 | _selectedValidData_T_97; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_113 = _selectedValidData_T_112 | _selectedValidData_T_98; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_114 = _selectedValidData_T_113 | _selectedValidData_T_99; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_115 = _selectedValidData_T_114 | _selectedValidData_T_100; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_116 = _selectedValidData_T_115 | _selectedValidData_T_101; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_117 = _selectedValidData_T_116 | _selectedValidData_T_102; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_118 = _selectedValidData_T_117 | _selectedValidData_T_103; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_119 = _selectedValidData_T_118 | _selectedValidData_T_104; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_120 = _selectedValidData_T_119 | _selectedValidData_T_105; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_121 = _selectedValidData_T_120 | _selectedValidData_T_106; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_122 = _selectedValidData_T_121 | _selectedValidData_T_107; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_3 = _selectedValidData_T_122 | _selectedValidData_T_108; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_124 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_125 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_126 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_127 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_128 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_129 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_130 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_131 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_132 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_133 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_134 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_135 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_136 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_137 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_138 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_139 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_140 = _selectedValidData_T_124 | _selectedValidData_T_125; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_141 = _selectedValidData_T_140 | _selectedValidData_T_126; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_142 = _selectedValidData_T_141 | _selectedValidData_T_127; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_143 = _selectedValidData_T_142 | _selectedValidData_T_128; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_144 = _selectedValidData_T_143 | _selectedValidData_T_129; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_145 = _selectedValidData_T_144 | _selectedValidData_T_130; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_146 = _selectedValidData_T_145 | _selectedValidData_T_131; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_147 = _selectedValidData_T_146 | _selectedValidData_T_132; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_148 = _selectedValidData_T_147 | _selectedValidData_T_133; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_149 = _selectedValidData_T_148 | _selectedValidData_T_134; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_150 = _selectedValidData_T_149 | _selectedValidData_T_135; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_151 = _selectedValidData_T_150 | _selectedValidData_T_136; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_152 = _selectedValidData_T_151 | _selectedValidData_T_137; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_153 = _selectedValidData_T_152 | _selectedValidData_T_138; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_4 = _selectedValidData_T_153 | _selectedValidData_T_139; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_155 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_156 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_157 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_158 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_159 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_160 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_161 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_162 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_163 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_164 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_165 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_166 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_167 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_168 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_169 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_170 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_171 = _selectedValidData_T_155 | _selectedValidData_T_156; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_172 = _selectedValidData_T_171 | _selectedValidData_T_157; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_173 = _selectedValidData_T_172 | _selectedValidData_T_158; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_174 = _selectedValidData_T_173 | _selectedValidData_T_159; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_175 = _selectedValidData_T_174 | _selectedValidData_T_160; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_176 = _selectedValidData_T_175 | _selectedValidData_T_161; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_177 = _selectedValidData_T_176 | _selectedValidData_T_162; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_178 = _selectedValidData_T_177 | _selectedValidData_T_163; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_179 = _selectedValidData_T_178 | _selectedValidData_T_164; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_180 = _selectedValidData_T_179 | _selectedValidData_T_165; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_181 = _selectedValidData_T_180 | _selectedValidData_T_166; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_182 = _selectedValidData_T_181 | _selectedValidData_T_167; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_183 = _selectedValidData_T_182 | _selectedValidData_T_168; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_184 = _selectedValidData_T_183 | _selectedValidData_T_169; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_5 = _selectedValidData_T_184 | _selectedValidData_T_170; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_186 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_187 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_188 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_189 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_190 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_191 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_192 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_193 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_194 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_195 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_196 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_197 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_198 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_199 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_200 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_201 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_202 = _selectedValidData_T_186 | _selectedValidData_T_187; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_203 = _selectedValidData_T_202 | _selectedValidData_T_188; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_204 = _selectedValidData_T_203 | _selectedValidData_T_189; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_205 = _selectedValidData_T_204 | _selectedValidData_T_190; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_206 = _selectedValidData_T_205 | _selectedValidData_T_191; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_207 = _selectedValidData_T_206 | _selectedValidData_T_192; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_208 = _selectedValidData_T_207 | _selectedValidData_T_193; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_209 = _selectedValidData_T_208 | _selectedValidData_T_194; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_210 = _selectedValidData_T_209 | _selectedValidData_T_195; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_211 = _selectedValidData_T_210 | _selectedValidData_T_196; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_212 = _selectedValidData_T_211 | _selectedValidData_T_197; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_213 = _selectedValidData_T_212 | _selectedValidData_T_198; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_214 = _selectedValidData_T_213 | _selectedValidData_T_199; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_215 = _selectedValidData_T_214 | _selectedValidData_T_200; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_6 = _selectedValidData_T_215 | _selectedValidData_T_201; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_217 = valid_tag_match_reg_0 ? forward_data_candidate_reg__0_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_218 = valid_tag_match_reg_1 ? forward_data_candidate_reg__1_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_219 = valid_tag_match_reg_2 ? forward_data_candidate_reg__2_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_220 = valid_tag_match_reg_3 ? forward_data_candidate_reg__3_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_221 = valid_tag_match_reg_4 ? forward_data_candidate_reg__4_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_222 = valid_tag_match_reg_5 ? forward_data_candidate_reg__5_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_223 = valid_tag_match_reg_6 ? forward_data_candidate_reg__6_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_224 = valid_tag_match_reg_7 ? forward_data_candidate_reg__7_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_225 = valid_tag_match_reg_8 ? forward_data_candidate_reg__8_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_226 = valid_tag_match_reg_9 ? forward_data_candidate_reg__9_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_227 = valid_tag_match_reg_10 ? forward_data_candidate_reg__10_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_228 = valid_tag_match_reg_11 ? forward_data_candidate_reg__11_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_229 = valid_tag_match_reg_12 ? forward_data_candidate_reg__12_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_230 = valid_tag_match_reg_13 ? forward_data_candidate_reg__13_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_231 = valid_tag_match_reg_14 ? forward_data_candidate_reg__14_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_232 = valid_tag_match_reg_15 ? forward_data_candidate_reg__15_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_233 = _selectedValidData_T_217 | _selectedValidData_T_218; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_234 = _selectedValidData_T_233 | _selectedValidData_T_219; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_235 = _selectedValidData_T_234 | _selectedValidData_T_220; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_236 = _selectedValidData_T_235 | _selectedValidData_T_221; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_237 = _selectedValidData_T_236 | _selectedValidData_T_222; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_238 = _selectedValidData_T_237 | _selectedValidData_T_223; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_239 = _selectedValidData_T_238 | _selectedValidData_T_224; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_240 = _selectedValidData_T_239 | _selectedValidData_T_225; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_241 = _selectedValidData_T_240 | _selectedValidData_T_226; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_242 = _selectedValidData_T_241 | _selectedValidData_T_227; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_243 = _selectedValidData_T_242 | _selectedValidData_T_228; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_244 = _selectedValidData_T_243 | _selectedValidData_T_229; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_245 = _selectedValidData_T_244 | _selectedValidData_T_230; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_246 = _selectedValidData_T_245 | _selectedValidData_T_231; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_0_7 = _selectedValidData_T_246 | _selectedValidData_T_232; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_15 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_0; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_0 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_0 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_0 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_0 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_0 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_0 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_0 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_0 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_0 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_0 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_0 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_0 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_0 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_0 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_0 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_0 |
    _selectedInflightMask_T_15; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_46 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_1; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_1 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_1 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_1 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_1 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_1 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_1 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_1 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_1 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_1 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_1 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_1 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_1 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_1 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_1 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_1 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_1 |
    _selectedInflightMask_T_46; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_77 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_2; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_2 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_2 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_2 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_2 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_2 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_2 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_2 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_2 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_2 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_2 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_2 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_2 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_2 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_2 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_2 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_2 |
    _selectedInflightMask_T_77; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_108 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_3; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_3 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_3 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_3 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_3 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_3 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_3 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_3 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_3 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_3 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_3 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_3 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_3 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_3 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_3 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_3 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_3 |
    _selectedInflightMask_T_108; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_139 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_4; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_4 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_4 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_4 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_4 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_4 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_4 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_4 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_4 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_4 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_4 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_4 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_4 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_4 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_4 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_4 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_4 |
    _selectedInflightMask_T_139; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_170 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_5; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_5 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_5 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_5 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_5 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_5 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_5 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_5 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_5 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_5 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_5 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_5 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_5 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_5 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_5 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_5 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_5 |
    _selectedInflightMask_T_170; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_201 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_6; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_6 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_6 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_6 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_6 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_6 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_6 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_6 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_6 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_6 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_6 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_6 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_6 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_6 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_6 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_6 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_6 |
    _selectedInflightMask_T_201; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_232 = inflight_tag_match_reg_15 & forward_mask_candidate_reg__15_7; // @[Mux.scala 27:73]
  wire  selectedInflightMask_0_7 = inflight_tag_match_reg_0 & forward_mask_candidate_reg__0_7 | inflight_tag_match_reg_1
     & forward_mask_candidate_reg__1_7 | inflight_tag_match_reg_2 & forward_mask_candidate_reg__2_7 |
    inflight_tag_match_reg_3 & forward_mask_candidate_reg__3_7 | inflight_tag_match_reg_4 &
    forward_mask_candidate_reg__4_7 | inflight_tag_match_reg_5 & forward_mask_candidate_reg__5_7 |
    inflight_tag_match_reg_6 & forward_mask_candidate_reg__6_7 | inflight_tag_match_reg_7 &
    forward_mask_candidate_reg__7_7 | inflight_tag_match_reg_8 & forward_mask_candidate_reg__8_7 |
    inflight_tag_match_reg_9 & forward_mask_candidate_reg__9_7 | inflight_tag_match_reg_10 &
    forward_mask_candidate_reg__10_7 | inflight_tag_match_reg_11 & forward_mask_candidate_reg__11_7 |
    inflight_tag_match_reg_12 & forward_mask_candidate_reg__12_7 | inflight_tag_match_reg_13 &
    forward_mask_candidate_reg__13_7 | inflight_tag_match_reg_14 & forward_mask_candidate_reg__14_7 |
    _selectedInflightMask_T_232; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_1 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_2 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_3 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_4 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_5 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_6 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_7 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_8 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_9 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_10 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_11 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_12 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_13 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_14 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_15 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_16 = _selectedInflightData_T | _selectedInflightData_T_1; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_17 = _selectedInflightData_T_16 | _selectedInflightData_T_2; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_18 = _selectedInflightData_T_17 | _selectedInflightData_T_3; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_19 = _selectedInflightData_T_18 | _selectedInflightData_T_4; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_20 = _selectedInflightData_T_19 | _selectedInflightData_T_5; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_21 = _selectedInflightData_T_20 | _selectedInflightData_T_6; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_22 = _selectedInflightData_T_21 | _selectedInflightData_T_7; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_23 = _selectedInflightData_T_22 | _selectedInflightData_T_8; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_24 = _selectedInflightData_T_23 | _selectedInflightData_T_9; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_25 = _selectedInflightData_T_24 | _selectedInflightData_T_10; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_26 = _selectedInflightData_T_25 | _selectedInflightData_T_11; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_27 = _selectedInflightData_T_26 | _selectedInflightData_T_12; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_28 = _selectedInflightData_T_27 | _selectedInflightData_T_13; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_29 = _selectedInflightData_T_28 | _selectedInflightData_T_14; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_0 = _selectedInflightData_T_29 | _selectedInflightData_T_15; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_31 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_32 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_33 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_34 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_35 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_36 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_37 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_38 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_39 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_40 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_41 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_42 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_43 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_44 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_45 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_46 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_47 = _selectedInflightData_T_31 | _selectedInflightData_T_32; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_48 = _selectedInflightData_T_47 | _selectedInflightData_T_33; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_49 = _selectedInflightData_T_48 | _selectedInflightData_T_34; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_50 = _selectedInflightData_T_49 | _selectedInflightData_T_35; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_51 = _selectedInflightData_T_50 | _selectedInflightData_T_36; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_52 = _selectedInflightData_T_51 | _selectedInflightData_T_37; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_53 = _selectedInflightData_T_52 | _selectedInflightData_T_38; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_54 = _selectedInflightData_T_53 | _selectedInflightData_T_39; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_55 = _selectedInflightData_T_54 | _selectedInflightData_T_40; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_56 = _selectedInflightData_T_55 | _selectedInflightData_T_41; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_57 = _selectedInflightData_T_56 | _selectedInflightData_T_42; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_58 = _selectedInflightData_T_57 | _selectedInflightData_T_43; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_59 = _selectedInflightData_T_58 | _selectedInflightData_T_44; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_60 = _selectedInflightData_T_59 | _selectedInflightData_T_45; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_1 = _selectedInflightData_T_60 | _selectedInflightData_T_46; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_62 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_63 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_64 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_65 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_66 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_67 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_68 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_69 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_70 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_71 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_72 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_73 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_74 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_75 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_76 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_77 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_78 = _selectedInflightData_T_62 | _selectedInflightData_T_63; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_79 = _selectedInflightData_T_78 | _selectedInflightData_T_64; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_80 = _selectedInflightData_T_79 | _selectedInflightData_T_65; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_81 = _selectedInflightData_T_80 | _selectedInflightData_T_66; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_82 = _selectedInflightData_T_81 | _selectedInflightData_T_67; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_83 = _selectedInflightData_T_82 | _selectedInflightData_T_68; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_84 = _selectedInflightData_T_83 | _selectedInflightData_T_69; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_85 = _selectedInflightData_T_84 | _selectedInflightData_T_70; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_86 = _selectedInflightData_T_85 | _selectedInflightData_T_71; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_87 = _selectedInflightData_T_86 | _selectedInflightData_T_72; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_88 = _selectedInflightData_T_87 | _selectedInflightData_T_73; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_89 = _selectedInflightData_T_88 | _selectedInflightData_T_74; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_90 = _selectedInflightData_T_89 | _selectedInflightData_T_75; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_91 = _selectedInflightData_T_90 | _selectedInflightData_T_76; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_2 = _selectedInflightData_T_91 | _selectedInflightData_T_77; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_93 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_94 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_95 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_96 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_97 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_98 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_99 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_100 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_101 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_102 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_103 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_104 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_105 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_106 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_107 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_108 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_109 = _selectedInflightData_T_93 | _selectedInflightData_T_94; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_110 = _selectedInflightData_T_109 | _selectedInflightData_T_95; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_111 = _selectedInflightData_T_110 | _selectedInflightData_T_96; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_112 = _selectedInflightData_T_111 | _selectedInflightData_T_97; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_113 = _selectedInflightData_T_112 | _selectedInflightData_T_98; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_114 = _selectedInflightData_T_113 | _selectedInflightData_T_99; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_115 = _selectedInflightData_T_114 | _selectedInflightData_T_100; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_116 = _selectedInflightData_T_115 | _selectedInflightData_T_101; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_117 = _selectedInflightData_T_116 | _selectedInflightData_T_102; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_118 = _selectedInflightData_T_117 | _selectedInflightData_T_103; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_119 = _selectedInflightData_T_118 | _selectedInflightData_T_104; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_120 = _selectedInflightData_T_119 | _selectedInflightData_T_105; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_121 = _selectedInflightData_T_120 | _selectedInflightData_T_106; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_122 = _selectedInflightData_T_121 | _selectedInflightData_T_107; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_3 = _selectedInflightData_T_122 | _selectedInflightData_T_108; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_124 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_125 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_126 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_127 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_128 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_129 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_130 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_131 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_132 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_133 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_134 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_135 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_136 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_137 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_138 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_139 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_140 = _selectedInflightData_T_124 | _selectedInflightData_T_125; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_141 = _selectedInflightData_T_140 | _selectedInflightData_T_126; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_142 = _selectedInflightData_T_141 | _selectedInflightData_T_127; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_143 = _selectedInflightData_T_142 | _selectedInflightData_T_128; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_144 = _selectedInflightData_T_143 | _selectedInflightData_T_129; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_145 = _selectedInflightData_T_144 | _selectedInflightData_T_130; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_146 = _selectedInflightData_T_145 | _selectedInflightData_T_131; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_147 = _selectedInflightData_T_146 | _selectedInflightData_T_132; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_148 = _selectedInflightData_T_147 | _selectedInflightData_T_133; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_149 = _selectedInflightData_T_148 | _selectedInflightData_T_134; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_150 = _selectedInflightData_T_149 | _selectedInflightData_T_135; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_151 = _selectedInflightData_T_150 | _selectedInflightData_T_136; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_152 = _selectedInflightData_T_151 | _selectedInflightData_T_137; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_153 = _selectedInflightData_T_152 | _selectedInflightData_T_138; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_4 = _selectedInflightData_T_153 | _selectedInflightData_T_139; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_155 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_156 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_157 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_158 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_159 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_160 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_161 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_162 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_163 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_164 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_165 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_166 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_167 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_168 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_169 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_170 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_171 = _selectedInflightData_T_155 | _selectedInflightData_T_156; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_172 = _selectedInflightData_T_171 | _selectedInflightData_T_157; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_173 = _selectedInflightData_T_172 | _selectedInflightData_T_158; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_174 = _selectedInflightData_T_173 | _selectedInflightData_T_159; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_175 = _selectedInflightData_T_174 | _selectedInflightData_T_160; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_176 = _selectedInflightData_T_175 | _selectedInflightData_T_161; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_177 = _selectedInflightData_T_176 | _selectedInflightData_T_162; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_178 = _selectedInflightData_T_177 | _selectedInflightData_T_163; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_179 = _selectedInflightData_T_178 | _selectedInflightData_T_164; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_180 = _selectedInflightData_T_179 | _selectedInflightData_T_165; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_181 = _selectedInflightData_T_180 | _selectedInflightData_T_166; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_182 = _selectedInflightData_T_181 | _selectedInflightData_T_167; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_183 = _selectedInflightData_T_182 | _selectedInflightData_T_168; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_184 = _selectedInflightData_T_183 | _selectedInflightData_T_169; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_5 = _selectedInflightData_T_184 | _selectedInflightData_T_170; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_186 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_187 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_188 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_189 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_190 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_191 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_192 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_193 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_194 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_195 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_196 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_197 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_198 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_199 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_200 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_201 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_202 = _selectedInflightData_T_186 | _selectedInflightData_T_187; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_203 = _selectedInflightData_T_202 | _selectedInflightData_T_188; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_204 = _selectedInflightData_T_203 | _selectedInflightData_T_189; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_205 = _selectedInflightData_T_204 | _selectedInflightData_T_190; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_206 = _selectedInflightData_T_205 | _selectedInflightData_T_191; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_207 = _selectedInflightData_T_206 | _selectedInflightData_T_192; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_208 = _selectedInflightData_T_207 | _selectedInflightData_T_193; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_209 = _selectedInflightData_T_208 | _selectedInflightData_T_194; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_210 = _selectedInflightData_T_209 | _selectedInflightData_T_195; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_211 = _selectedInflightData_T_210 | _selectedInflightData_T_196; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_212 = _selectedInflightData_T_211 | _selectedInflightData_T_197; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_213 = _selectedInflightData_T_212 | _selectedInflightData_T_198; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_214 = _selectedInflightData_T_213 | _selectedInflightData_T_199; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_215 = _selectedInflightData_T_214 | _selectedInflightData_T_200; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_6 = _selectedInflightData_T_215 | _selectedInflightData_T_201; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_217 = inflight_tag_match_reg_0 ? forward_data_candidate_reg__0_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_218 = inflight_tag_match_reg_1 ? forward_data_candidate_reg__1_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_219 = inflight_tag_match_reg_2 ? forward_data_candidate_reg__2_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_220 = inflight_tag_match_reg_3 ? forward_data_candidate_reg__3_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_221 = inflight_tag_match_reg_4 ? forward_data_candidate_reg__4_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_222 = inflight_tag_match_reg_5 ? forward_data_candidate_reg__5_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_223 = inflight_tag_match_reg_6 ? forward_data_candidate_reg__6_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_224 = inflight_tag_match_reg_7 ? forward_data_candidate_reg__7_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_225 = inflight_tag_match_reg_8 ? forward_data_candidate_reg__8_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_226 = inflight_tag_match_reg_9 ? forward_data_candidate_reg__9_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_227 = inflight_tag_match_reg_10 ? forward_data_candidate_reg__10_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_228 = inflight_tag_match_reg_11 ? forward_data_candidate_reg__11_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_229 = inflight_tag_match_reg_12 ? forward_data_candidate_reg__12_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_230 = inflight_tag_match_reg_13 ? forward_data_candidate_reg__13_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_231 = inflight_tag_match_reg_14 ? forward_data_candidate_reg__14_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_232 = inflight_tag_match_reg_15 ? forward_data_candidate_reg__15_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_233 = _selectedInflightData_T_217 | _selectedInflightData_T_218; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_234 = _selectedInflightData_T_233 | _selectedInflightData_T_219; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_235 = _selectedInflightData_T_234 | _selectedInflightData_T_220; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_236 = _selectedInflightData_T_235 | _selectedInflightData_T_221; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_237 = _selectedInflightData_T_236 | _selectedInflightData_T_222; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_238 = _selectedInflightData_T_237 | _selectedInflightData_T_223; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_239 = _selectedInflightData_T_238 | _selectedInflightData_T_224; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_240 = _selectedInflightData_T_239 | _selectedInflightData_T_225; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_241 = _selectedInflightData_T_240 | _selectedInflightData_T_226; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_242 = _selectedInflightData_T_241 | _selectedInflightData_T_227; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_243 = _selectedInflightData_T_242 | _selectedInflightData_T_228; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_244 = _selectedInflightData_T_243 | _selectedInflightData_T_229; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_245 = _selectedInflightData_T_244 | _selectedInflightData_T_230; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_246 = _selectedInflightData_T_245 | _selectedInflightData_T_231; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_0_7 = _selectedInflightData_T_246 | _selectedInflightData_T_232; // @[Mux.scala 27:73]
  wire  vtag_matches_1_0 = vtag_0 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_1 = vtag_1 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_2 = vtag_2 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_3 = vtag_3 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_4 = vtag_4 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_5 = vtag_5 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_6 = vtag_6 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_7 = vtag_7 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_8 = vtag_8 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_9 = vtag_9 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_10 = vtag_10 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_11 = vtag_11 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_12 = vtag_12 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_13 = vtag_13 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_14 = vtag_14 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  wire  vtag_matches_1_15 = vtag_15 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
  reg  valid_tag_match_reg_0_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_1_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_2_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_3_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_4_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_5_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_6_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_7_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_8_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_9_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_10_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_11_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_12_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_13_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_14_1; // @[Sbuffer.scala 816:60]
  reg  valid_tag_match_reg_15_1; // @[Sbuffer.scala 816:60]
  reg  inflight_tag_match_reg_0_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_1_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_2_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_3_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_4_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_5_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_6_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_7_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_8_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_9_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_10_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_11_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_12_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_13_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_14_1; // @[Sbuffer.scala 817:66]
  reg  inflight_tag_match_reg_15_1; // @[Sbuffer.scala 817:66]
  wire  _GEN_5663 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_0 : _GEN_1948; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5664 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_0 : _GEN_5663; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5665 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_0 : _GEN_5664; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5666 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_0 : _GEN_5665; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5671 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_1 : _GEN_1932; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5672 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_1 : _GEN_5671; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5673 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_1 : _GEN_5672; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5674 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_1 : _GEN_5673; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5679 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_2 : _GEN_1980; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5680 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_2 : _GEN_5679; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5681 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_2 : _GEN_5680; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5682 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_2 : _GEN_5681; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5687 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_3 : _GEN_1964; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5688 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_3 : _GEN_5687; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5689 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_3 : _GEN_5688; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5690 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_3 : _GEN_5689; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5695 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_4 : _GEN_2012; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5696 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_4 : _GEN_5695; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5697 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_4 : _GEN_5696; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5698 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_4 : _GEN_5697; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5703 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_5 : _GEN_1996; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5704 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_5 : _GEN_5703; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5705 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_5 : _GEN_5704; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5706 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_5 : _GEN_5705; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5711 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_6 : _GEN_2044; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5712 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_6 : _GEN_5711; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5713 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_6 : _GEN_5712; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5714 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_6 : _GEN_5713; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5719 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_1_7 : _GEN_2028; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5720 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_2_7 : _GEN_5719; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5721 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_3_7 : _GEN_5720; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5722 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_0_4_7 : _GEN_5721; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5727 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_0 : dataModule_io_maskOut_1_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5728 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_0 : _GEN_5727; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5729 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_0 : _GEN_5728; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5730 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_0 : _GEN_5729; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5735 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_1 : dataModule_io_maskOut_1_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5736 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_1 : _GEN_5735; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5737 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_1 : _GEN_5736; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5738 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_1 : _GEN_5737; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5743 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_2 : dataModule_io_maskOut_1_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5744 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_2 : _GEN_5743; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5745 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_2 : _GEN_5744; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5746 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_2 : _GEN_5745; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5751 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_3 : dataModule_io_maskOut_1_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5752 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_3 : _GEN_5751; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5753 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_3 : _GEN_5752; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5754 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_3 : _GEN_5753; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5759 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_4 : dataModule_io_maskOut_1_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5760 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_4 : _GEN_5759; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5761 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_4 : _GEN_5760; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5762 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_4 : _GEN_5761; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5767 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_5 : dataModule_io_maskOut_1_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5768 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_5 : _GEN_5767; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5769 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_5 : _GEN_5768; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5770 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_5 : _GEN_5769; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5775 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_6 : dataModule_io_maskOut_1_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5776 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_6 : _GEN_5775; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5777 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_6 : _GEN_5776; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5778 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_6 : _GEN_5777; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5783 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_1_7 : dataModule_io_maskOut_1_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5784 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_2_7 : _GEN_5783; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5785 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_3_7 : _GEN_5784; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5786 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_1_4_7 : _GEN_5785; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5791 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_0 : dataModule_io_maskOut_2_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5792 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_0 : _GEN_5791; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5793 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_0 : _GEN_5792; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5794 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_0 : _GEN_5793; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5799 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_1 : dataModule_io_maskOut_2_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5800 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_1 : _GEN_5799; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5801 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_1 : _GEN_5800; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5802 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_1 : _GEN_5801; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5807 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_2 : dataModule_io_maskOut_2_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5808 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_2 : _GEN_5807; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5809 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_2 : _GEN_5808; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5810 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_2 : _GEN_5809; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5815 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_3 : dataModule_io_maskOut_2_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5816 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_3 : _GEN_5815; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5817 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_3 : _GEN_5816; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5818 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_3 : _GEN_5817; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5823 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_4 : dataModule_io_maskOut_2_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5824 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_4 : _GEN_5823; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5825 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_4 : _GEN_5824; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5826 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_4 : _GEN_5825; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5831 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_5 : dataModule_io_maskOut_2_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5832 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_5 : _GEN_5831; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5833 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_5 : _GEN_5832; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5834 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_5 : _GEN_5833; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5839 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_6 : dataModule_io_maskOut_2_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5840 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_6 : _GEN_5839; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5841 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_6 : _GEN_5840; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5842 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_6 : _GEN_5841; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5847 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_1_7 : dataModule_io_maskOut_2_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5848 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_2_7 : _GEN_5847; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5849 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_3_7 : _GEN_5848; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5850 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_2_4_7 : _GEN_5849; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5855 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_0 : dataModule_io_maskOut_3_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5856 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_0 : _GEN_5855; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5857 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_0 : _GEN_5856; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5858 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_0 : _GEN_5857; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5863 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_1 : dataModule_io_maskOut_3_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5864 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_1 : _GEN_5863; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5865 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_1 : _GEN_5864; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5866 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_1 : _GEN_5865; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5871 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_2 : dataModule_io_maskOut_3_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5872 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_2 : _GEN_5871; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5873 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_2 : _GEN_5872; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5874 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_2 : _GEN_5873; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5879 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_3 : dataModule_io_maskOut_3_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5880 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_3 : _GEN_5879; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5881 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_3 : _GEN_5880; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5882 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_3 : _GEN_5881; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5887 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_4 : dataModule_io_maskOut_3_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5888 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_4 : _GEN_5887; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5889 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_4 : _GEN_5888; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5890 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_4 : _GEN_5889; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5895 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_5 : dataModule_io_maskOut_3_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5896 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_5 : _GEN_5895; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5897 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_5 : _GEN_5896; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5898 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_5 : _GEN_5897; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5903 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_6 : dataModule_io_maskOut_3_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5904 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_6 : _GEN_5903; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5905 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_6 : _GEN_5904; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5906 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_6 : _GEN_5905; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5911 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_1_7 : dataModule_io_maskOut_3_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5912 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_2_7 : _GEN_5911; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5913 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_3_7 : _GEN_5912; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5914 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_3_4_7 : _GEN_5913; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5919 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_0 : dataModule_io_maskOut_4_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5920 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_0 : _GEN_5919; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5921 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_0 : _GEN_5920; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5922 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_0 : _GEN_5921; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5927 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_1 : dataModule_io_maskOut_4_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5928 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_1 : _GEN_5927; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5929 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_1 : _GEN_5928; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5930 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_1 : _GEN_5929; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5935 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_2 : dataModule_io_maskOut_4_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5936 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_2 : _GEN_5935; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5937 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_2 : _GEN_5936; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5938 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_2 : _GEN_5937; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5943 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_3 : dataModule_io_maskOut_4_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5944 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_3 : _GEN_5943; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5945 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_3 : _GEN_5944; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5946 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_3 : _GEN_5945; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5951 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_4 : dataModule_io_maskOut_4_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5952 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_4 : _GEN_5951; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5953 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_4 : _GEN_5952; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5954 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_4 : _GEN_5953; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5959 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_5 : dataModule_io_maskOut_4_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5960 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_5 : _GEN_5959; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5961 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_5 : _GEN_5960; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5962 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_5 : _GEN_5961; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5967 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_6 : dataModule_io_maskOut_4_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5968 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_6 : _GEN_5967; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5969 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_6 : _GEN_5968; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5970 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_6 : _GEN_5969; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5975 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_1_7 : dataModule_io_maskOut_4_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5976 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_2_7 : _GEN_5975; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5977 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_3_7 : _GEN_5976; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5978 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_4_4_7 : _GEN_5977; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5983 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_0 : dataModule_io_maskOut_5_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5984 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_0 : _GEN_5983; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5985 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_0 : _GEN_5984; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5986 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_0 : _GEN_5985; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5991 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_1 : dataModule_io_maskOut_5_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5992 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_1 : _GEN_5991; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5993 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_1 : _GEN_5992; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5994 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_1 : _GEN_5993; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_5999 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_2 : dataModule_io_maskOut_5_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6000 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_2 : _GEN_5999; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6001 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_2 : _GEN_6000; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6002 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_2 : _GEN_6001; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6007 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_3 : dataModule_io_maskOut_5_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6008 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_3 : _GEN_6007; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6009 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_3 : _GEN_6008; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6010 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_3 : _GEN_6009; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6015 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_4 : dataModule_io_maskOut_5_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6016 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_4 : _GEN_6015; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6017 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_4 : _GEN_6016; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6018 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_4 : _GEN_6017; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6023 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_5 : dataModule_io_maskOut_5_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6024 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_5 : _GEN_6023; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6025 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_5 : _GEN_6024; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6026 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_5 : _GEN_6025; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6031 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_6 : dataModule_io_maskOut_5_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6032 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_6 : _GEN_6031; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6033 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_6 : _GEN_6032; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6034 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_6 : _GEN_6033; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6039 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_1_7 : dataModule_io_maskOut_5_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6040 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_2_7 : _GEN_6039; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6041 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_3_7 : _GEN_6040; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6042 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_5_4_7 : _GEN_6041; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6047 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_0 : dataModule_io_maskOut_6_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6048 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_0 : _GEN_6047; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6049 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_0 : _GEN_6048; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6050 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_0 : _GEN_6049; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6055 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_1 : dataModule_io_maskOut_6_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6056 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_1 : _GEN_6055; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6057 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_1 : _GEN_6056; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6058 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_1 : _GEN_6057; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6063 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_2 : dataModule_io_maskOut_6_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6064 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_2 : _GEN_6063; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6065 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_2 : _GEN_6064; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6066 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_2 : _GEN_6065; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6071 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_3 : dataModule_io_maskOut_6_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6072 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_3 : _GEN_6071; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6073 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_3 : _GEN_6072; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6074 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_3 : _GEN_6073; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6079 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_4 : dataModule_io_maskOut_6_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6080 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_4 : _GEN_6079; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6081 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_4 : _GEN_6080; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6082 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_4 : _GEN_6081; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6087 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_5 : dataModule_io_maskOut_6_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6088 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_5 : _GEN_6087; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6089 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_5 : _GEN_6088; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6090 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_5 : _GEN_6089; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6095 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_6 : dataModule_io_maskOut_6_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6096 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_6 : _GEN_6095; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6097 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_6 : _GEN_6096; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6098 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_6 : _GEN_6097; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6103 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_1_7 : dataModule_io_maskOut_6_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6104 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_2_7 : _GEN_6103; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6105 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_3_7 : _GEN_6104; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6106 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_6_4_7 : _GEN_6105; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6111 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_0 : dataModule_io_maskOut_7_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6112 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_0 : _GEN_6111; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6113 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_0 : _GEN_6112; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6114 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_0 : _GEN_6113; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6119 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_1 : dataModule_io_maskOut_7_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6120 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_1 : _GEN_6119; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6121 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_1 : _GEN_6120; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6122 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_1 : _GEN_6121; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6127 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_2 : dataModule_io_maskOut_7_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6128 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_2 : _GEN_6127; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6129 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_2 : _GEN_6128; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6130 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_2 : _GEN_6129; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6135 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_3 : dataModule_io_maskOut_7_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6136 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_3 : _GEN_6135; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6137 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_3 : _GEN_6136; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6138 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_3 : _GEN_6137; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6143 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_4 : dataModule_io_maskOut_7_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6144 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_4 : _GEN_6143; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6145 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_4 : _GEN_6144; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6146 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_4 : _GEN_6145; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6151 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_5 : dataModule_io_maskOut_7_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6152 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_5 : _GEN_6151; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6153 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_5 : _GEN_6152; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6154 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_5 : _GEN_6153; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6159 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_6 : dataModule_io_maskOut_7_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6160 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_6 : _GEN_6159; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6161 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_6 : _GEN_6160; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6162 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_6 : _GEN_6161; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6167 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_1_7 : dataModule_io_maskOut_7_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6168 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_2_7 : _GEN_6167; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6169 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_3_7 : _GEN_6168; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6170 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_7_4_7 : _GEN_6169; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6175 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_0 : dataModule_io_maskOut_8_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6176 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_0 : _GEN_6175; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6177 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_0 : _GEN_6176; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6178 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_0 : _GEN_6177; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6183 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_1 : dataModule_io_maskOut_8_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6184 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_1 : _GEN_6183; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6185 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_1 : _GEN_6184; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6186 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_1 : _GEN_6185; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6191 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_2 : dataModule_io_maskOut_8_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6192 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_2 : _GEN_6191; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6193 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_2 : _GEN_6192; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6194 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_2 : _GEN_6193; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6199 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_3 : dataModule_io_maskOut_8_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6200 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_3 : _GEN_6199; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6201 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_3 : _GEN_6200; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6202 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_3 : _GEN_6201; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6207 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_4 : dataModule_io_maskOut_8_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6208 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_4 : _GEN_6207; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6209 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_4 : _GEN_6208; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6210 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_4 : _GEN_6209; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6215 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_5 : dataModule_io_maskOut_8_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6216 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_5 : _GEN_6215; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6217 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_5 : _GEN_6216; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6218 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_5 : _GEN_6217; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6223 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_6 : dataModule_io_maskOut_8_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6224 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_6 : _GEN_6223; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6225 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_6 : _GEN_6224; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6226 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_6 : _GEN_6225; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6231 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_1_7 : dataModule_io_maskOut_8_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6232 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_2_7 : _GEN_6231; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6233 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_3_7 : _GEN_6232; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6234 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_8_4_7 : _GEN_6233; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6239 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_0 : dataModule_io_maskOut_9_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6240 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_0 : _GEN_6239; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6241 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_0 : _GEN_6240; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6242 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_0 : _GEN_6241; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6247 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_1 : dataModule_io_maskOut_9_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6248 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_1 : _GEN_6247; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6249 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_1 : _GEN_6248; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6250 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_1 : _GEN_6249; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6255 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_2 : dataModule_io_maskOut_9_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6256 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_2 : _GEN_6255; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6257 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_2 : _GEN_6256; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6258 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_2 : _GEN_6257; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6263 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_3 : dataModule_io_maskOut_9_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6264 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_3 : _GEN_6263; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6265 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_3 : _GEN_6264; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6266 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_3 : _GEN_6265; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6271 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_4 : dataModule_io_maskOut_9_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6272 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_4 : _GEN_6271; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6273 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_4 : _GEN_6272; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6274 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_4 : _GEN_6273; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6279 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_5 : dataModule_io_maskOut_9_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6280 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_5 : _GEN_6279; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6281 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_5 : _GEN_6280; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6282 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_5 : _GEN_6281; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6287 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_6 : dataModule_io_maskOut_9_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6288 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_6 : _GEN_6287; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6289 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_6 : _GEN_6288; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6290 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_6 : _GEN_6289; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6295 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_1_7 : dataModule_io_maskOut_9_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6296 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_2_7 : _GEN_6295; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6297 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_3_7 : _GEN_6296; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6298 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_9_4_7 : _GEN_6297; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6303 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_0 : dataModule_io_maskOut_10_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6304 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_0 : _GEN_6303; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6305 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_0 : _GEN_6304; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6306 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_0 : _GEN_6305; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6311 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_1 : dataModule_io_maskOut_10_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6312 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_1 : _GEN_6311; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6313 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_1 : _GEN_6312; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6314 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_1 : _GEN_6313; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6319 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_2 : dataModule_io_maskOut_10_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6320 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_2 : _GEN_6319; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6321 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_2 : _GEN_6320; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6322 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_2 : _GEN_6321; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6327 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_3 : dataModule_io_maskOut_10_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6328 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_3 : _GEN_6327; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6329 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_3 : _GEN_6328; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6330 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_3 : _GEN_6329; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6335 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_4 : dataModule_io_maskOut_10_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6336 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_4 : _GEN_6335; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6337 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_4 : _GEN_6336; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6338 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_4 : _GEN_6337; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6343 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_5 : dataModule_io_maskOut_10_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6344 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_5 : _GEN_6343; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6345 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_5 : _GEN_6344; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6346 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_5 : _GEN_6345; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6351 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_6 : dataModule_io_maskOut_10_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6352 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_6 : _GEN_6351; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6353 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_6 : _GEN_6352; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6354 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_6 : _GEN_6353; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6359 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_1_7 : dataModule_io_maskOut_10_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6360 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_2_7 : _GEN_6359; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6361 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_3_7 : _GEN_6360; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6362 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_10_4_7 : _GEN_6361; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6367 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_0 : dataModule_io_maskOut_11_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6368 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_0 : _GEN_6367; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6369 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_0 : _GEN_6368; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6370 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_0 : _GEN_6369; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6375 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_1 : dataModule_io_maskOut_11_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6376 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_1 : _GEN_6375; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6377 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_1 : _GEN_6376; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6378 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_1 : _GEN_6377; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6383 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_2 : dataModule_io_maskOut_11_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6384 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_2 : _GEN_6383; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6385 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_2 : _GEN_6384; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6386 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_2 : _GEN_6385; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6391 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_3 : dataModule_io_maskOut_11_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6392 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_3 : _GEN_6391; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6393 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_3 : _GEN_6392; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6394 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_3 : _GEN_6393; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6399 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_4 : dataModule_io_maskOut_11_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6400 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_4 : _GEN_6399; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6401 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_4 : _GEN_6400; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6402 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_4 : _GEN_6401; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6407 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_5 : dataModule_io_maskOut_11_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6408 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_5 : _GEN_6407; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6409 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_5 : _GEN_6408; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6410 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_5 : _GEN_6409; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6415 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_6 : dataModule_io_maskOut_11_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6416 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_6 : _GEN_6415; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6417 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_6 : _GEN_6416; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6418 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_6 : _GEN_6417; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6423 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_1_7 : dataModule_io_maskOut_11_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6424 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_2_7 : _GEN_6423; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6425 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_3_7 : _GEN_6424; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6426 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_11_4_7 : _GEN_6425; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6431 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_0 : dataModule_io_maskOut_12_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6432 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_0 : _GEN_6431; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6433 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_0 : _GEN_6432; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6434 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_0 : _GEN_6433; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6439 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_1 : dataModule_io_maskOut_12_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6440 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_1 : _GEN_6439; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6441 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_1 : _GEN_6440; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6442 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_1 : _GEN_6441; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6447 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_2 : dataModule_io_maskOut_12_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6448 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_2 : _GEN_6447; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6449 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_2 : _GEN_6448; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6450 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_2 : _GEN_6449; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6455 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_3 : dataModule_io_maskOut_12_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6456 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_3 : _GEN_6455; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6457 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_3 : _GEN_6456; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6458 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_3 : _GEN_6457; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6463 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_4 : dataModule_io_maskOut_12_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6464 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_4 : _GEN_6463; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6465 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_4 : _GEN_6464; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6466 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_4 : _GEN_6465; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6471 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_5 : dataModule_io_maskOut_12_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6472 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_5 : _GEN_6471; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6473 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_5 : _GEN_6472; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6474 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_5 : _GEN_6473; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6479 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_6 : dataModule_io_maskOut_12_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6480 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_6 : _GEN_6479; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6481 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_6 : _GEN_6480; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6482 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_6 : _GEN_6481; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6487 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_1_7 : dataModule_io_maskOut_12_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6488 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_2_7 : _GEN_6487; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6489 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_3_7 : _GEN_6488; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6490 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_12_4_7 : _GEN_6489; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6495 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_0 : dataModule_io_maskOut_13_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6496 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_0 : _GEN_6495; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6497 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_0 : _GEN_6496; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6498 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_0 : _GEN_6497; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6503 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_1 : dataModule_io_maskOut_13_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6504 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_1 : _GEN_6503; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6505 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_1 : _GEN_6504; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6506 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_1 : _GEN_6505; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6511 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_2 : dataModule_io_maskOut_13_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6512 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_2 : _GEN_6511; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6513 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_2 : _GEN_6512; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6514 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_2 : _GEN_6513; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6519 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_3 : dataModule_io_maskOut_13_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6520 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_3 : _GEN_6519; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6521 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_3 : _GEN_6520; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6522 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_3 : _GEN_6521; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6527 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_4 : dataModule_io_maskOut_13_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6528 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_4 : _GEN_6527; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6529 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_4 : _GEN_6528; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6530 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_4 : _GEN_6529; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6535 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_5 : dataModule_io_maskOut_13_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6536 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_5 : _GEN_6535; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6537 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_5 : _GEN_6536; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6538 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_5 : _GEN_6537; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6543 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_6 : dataModule_io_maskOut_13_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6544 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_6 : _GEN_6543; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6545 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_6 : _GEN_6544; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6546 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_6 : _GEN_6545; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6551 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_1_7 : dataModule_io_maskOut_13_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6552 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_2_7 : _GEN_6551; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6553 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_3_7 : _GEN_6552; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6554 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_13_4_7 : _GEN_6553; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6559 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_0 : dataModule_io_maskOut_14_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6560 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_0 : _GEN_6559; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6561 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_0 : _GEN_6560; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6562 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_0 : _GEN_6561; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6567 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_1 : dataModule_io_maskOut_14_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6568 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_1 : _GEN_6567; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6569 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_1 : _GEN_6568; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6570 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_1 : _GEN_6569; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6575 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_2 : dataModule_io_maskOut_14_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6576 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_2 : _GEN_6575; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6577 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_2 : _GEN_6576; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6578 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_2 : _GEN_6577; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6583 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_3 : dataModule_io_maskOut_14_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6584 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_3 : _GEN_6583; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6585 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_3 : _GEN_6584; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6586 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_3 : _GEN_6585; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6591 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_4 : dataModule_io_maskOut_14_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6592 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_4 : _GEN_6591; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6593 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_4 : _GEN_6592; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6594 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_4 : _GEN_6593; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6599 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_5 : dataModule_io_maskOut_14_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6600 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_5 : _GEN_6599; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6601 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_5 : _GEN_6600; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6602 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_5 : _GEN_6601; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6607 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_6 : dataModule_io_maskOut_14_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6608 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_6 : _GEN_6607; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6609 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_6 : _GEN_6608; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6610 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_6 : _GEN_6609; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6615 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_1_7 : dataModule_io_maskOut_14_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6616 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_2_7 : _GEN_6615; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6617 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_3_7 : _GEN_6616; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6618 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_14_4_7 : _GEN_6617; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6623 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_0 : dataModule_io_maskOut_15_0_0; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6624 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_0 : _GEN_6623; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6625 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_0 : _GEN_6624; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6626 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_0 : _GEN_6625; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6631 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_1 : dataModule_io_maskOut_15_0_1; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6632 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_1 : _GEN_6631; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6633 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_1 : _GEN_6632; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6634 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_1 : _GEN_6633; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6639 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_2 : dataModule_io_maskOut_15_0_2; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6640 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_2 : _GEN_6639; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6641 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_2 : _GEN_6640; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6642 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_2 : _GEN_6641; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6647 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_3 : dataModule_io_maskOut_15_0_3; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6648 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_3 : _GEN_6647; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6649 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_3 : _GEN_6648; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6650 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_3 : _GEN_6649; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6655 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_4 : dataModule_io_maskOut_15_0_4; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6656 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_4 : _GEN_6655; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6657 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_4 : _GEN_6656; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6658 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_4 : _GEN_6657; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6663 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_5 : dataModule_io_maskOut_15_0_5; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6664 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_5 : _GEN_6663; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6665 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_5 : _GEN_6664; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6666 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_5 : _GEN_6665; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6671 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_6 : dataModule_io_maskOut_15_0_6; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6672 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_6 : _GEN_6671; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6673 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_6 : _GEN_6672; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6674 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_6 : _GEN_6673; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6679 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_1_7 : dataModule_io_maskOut_15_0_7; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6680 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_2_7 : _GEN_6679; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6681 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_3_7 : _GEN_6680; // @[Sbuffer.scala 820:{14,14}]
  wire  _GEN_6682 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_maskOut_15_4_7 : _GEN_6681; // @[Sbuffer.scala 820:{14,14}]
  reg  forward_mask_candidate_reg_1_0_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_0_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_1_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_2_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_3_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_4_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_5_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_6_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_7_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_8_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_9_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_10_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_11_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_12_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_13_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_14_7; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_0; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_1; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_2; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_3; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_4; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_5; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_6; // @[Reg.scala 19:16]
  reg  forward_mask_candidate_reg_1_15_7; // @[Reg.scala 19:16]
  wire [7:0] _GEN_6815 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_0 : _GEN_924; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6816 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_0 : _GEN_6815; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6817 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_0 : _GEN_6816; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6818 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_0 : _GEN_6817; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6823 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_1 : _GEN_908; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6824 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_1 : _GEN_6823; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6825 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_1 : _GEN_6824; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6826 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_1 : _GEN_6825; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6831 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_2 : _GEN_956; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6832 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_2 : _GEN_6831; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6833 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_2 : _GEN_6832; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6834 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_2 : _GEN_6833; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6839 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_3 : _GEN_940; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6840 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_3 : _GEN_6839; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6841 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_3 : _GEN_6840; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6842 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_3 : _GEN_6841; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6847 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_4 : _GEN_988; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6848 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_4 : _GEN_6847; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6849 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_4 : _GEN_6848; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6850 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_4 : _GEN_6849; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6855 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_5 : _GEN_972; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6856 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_5 : _GEN_6855; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6857 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_5 : _GEN_6856; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6858 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_5 : _GEN_6857; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6863 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_6 : _GEN_1020; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6864 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_6 : _GEN_6863; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6865 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_6 : _GEN_6864; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6866 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_6 : _GEN_6865; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6871 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_1_7 : _GEN_1004; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6872 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_2_7 : _GEN_6871; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6873 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_3_7 : _GEN_6872; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6874 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_0_4_7 : _GEN_6873; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6879 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_0 : _GEN_4509; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6880 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_0 : _GEN_6879; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6881 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_0 : _GEN_6880; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6882 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_0 : _GEN_6881; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6887 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_1 : _GEN_4517; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6888 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_1 : _GEN_6887; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6889 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_1 : _GEN_6888; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6890 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_1 : _GEN_6889; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6895 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_2 : _GEN_4525; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6896 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_2 : _GEN_6895; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6897 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_2 : _GEN_6896; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6898 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_2 : _GEN_6897; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6903 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_3 : _GEN_4533; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6904 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_3 : _GEN_6903; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6905 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_3 : _GEN_6904; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6906 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_3 : _GEN_6905; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6911 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_4 : _GEN_4541; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6912 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_4 : _GEN_6911; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6913 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_4 : _GEN_6912; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6914 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_4 : _GEN_6913; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6919 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_5 : _GEN_4549; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6920 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_5 : _GEN_6919; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6921 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_5 : _GEN_6920; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6922 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_5 : _GEN_6921; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6927 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_6 : _GEN_4557; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6928 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_6 : _GEN_6927; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6929 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_6 : _GEN_6928; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6930 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_6 : _GEN_6929; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6935 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_1_7 : _GEN_4565; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6936 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_2_7 : _GEN_6935; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6937 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_3_7 : _GEN_6936; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6938 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_1_4_7 : _GEN_6937; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6943 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_0 : _GEN_4573; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6944 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_0 : _GEN_6943; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6945 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_0 : _GEN_6944; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6946 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_0 : _GEN_6945; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6951 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_1 : _GEN_4581; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6952 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_1 : _GEN_6951; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6953 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_1 : _GEN_6952; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6954 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_1 : _GEN_6953; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6959 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_2 : _GEN_4589; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6960 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_2 : _GEN_6959; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6961 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_2 : _GEN_6960; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6962 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_2 : _GEN_6961; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6967 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_3 : _GEN_4597; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6968 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_3 : _GEN_6967; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6969 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_3 : _GEN_6968; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6970 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_3 : _GEN_6969; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6975 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_4 : _GEN_4605; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6976 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_4 : _GEN_6975; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6977 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_4 : _GEN_6976; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6978 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_4 : _GEN_6977; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6983 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_5 : _GEN_4613; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6984 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_5 : _GEN_6983; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6985 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_5 : _GEN_6984; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6986 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_5 : _GEN_6985; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6991 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_6 : _GEN_4621; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6992 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_6 : _GEN_6991; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6993 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_6 : _GEN_6992; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6994 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_6 : _GEN_6993; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_6999 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_1_7 : _GEN_4629; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7000 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_2_7 : _GEN_6999; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7001 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_3_7 : _GEN_7000; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7002 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_2_4_7 : _GEN_7001; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7007 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_0 : _GEN_4637; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7008 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_0 : _GEN_7007; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7009 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_0 : _GEN_7008; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7010 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_0 : _GEN_7009; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7015 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_1 : _GEN_4645; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7016 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_1 : _GEN_7015; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7017 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_1 : _GEN_7016; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7018 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_1 : _GEN_7017; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7023 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_2 : _GEN_4653; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7024 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_2 : _GEN_7023; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7025 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_2 : _GEN_7024; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7026 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_2 : _GEN_7025; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7031 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_3 : _GEN_4661; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7032 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_3 : _GEN_7031; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7033 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_3 : _GEN_7032; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7034 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_3 : _GEN_7033; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7039 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_4 : _GEN_4669; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7040 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_4 : _GEN_7039; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7041 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_4 : _GEN_7040; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7042 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_4 : _GEN_7041; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7047 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_5 : _GEN_4677; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7048 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_5 : _GEN_7047; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7049 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_5 : _GEN_7048; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7050 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_5 : _GEN_7049; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7055 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_6 : _GEN_4685; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7056 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_6 : _GEN_7055; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7057 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_6 : _GEN_7056; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7058 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_6 : _GEN_7057; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7063 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_1_7 : _GEN_4693; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7064 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_2_7 : _GEN_7063; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7065 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_3_7 : _GEN_7064; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7066 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_3_4_7 : _GEN_7065; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7071 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_0 : _GEN_4701; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7072 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_0 : _GEN_7071; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7073 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_0 : _GEN_7072; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7074 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_0 : _GEN_7073; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7079 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_1 : _GEN_4709; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7080 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_1 : _GEN_7079; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7081 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_1 : _GEN_7080; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7082 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_1 : _GEN_7081; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7087 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_2 : _GEN_4717; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7088 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_2 : _GEN_7087; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7089 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_2 : _GEN_7088; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7090 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_2 : _GEN_7089; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7095 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_3 : _GEN_4725; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7096 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_3 : _GEN_7095; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7097 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_3 : _GEN_7096; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7098 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_3 : _GEN_7097; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7103 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_4 : _GEN_4733; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7104 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_4 : _GEN_7103; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7105 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_4 : _GEN_7104; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7106 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_4 : _GEN_7105; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7111 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_5 : _GEN_4741; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7112 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_5 : _GEN_7111; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7113 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_5 : _GEN_7112; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7114 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_5 : _GEN_7113; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7119 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_6 : _GEN_4749; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7120 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_6 : _GEN_7119; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7121 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_6 : _GEN_7120; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7122 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_6 : _GEN_7121; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7127 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_1_7 : _GEN_4757; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7128 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_2_7 : _GEN_7127; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7129 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_3_7 : _GEN_7128; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7130 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_4_4_7 : _GEN_7129; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7135 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_0 : _GEN_4765; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7136 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_0 : _GEN_7135; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7137 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_0 : _GEN_7136; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7138 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_0 : _GEN_7137; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7143 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_1 : _GEN_4773; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7144 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_1 : _GEN_7143; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7145 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_1 : _GEN_7144; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7146 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_1 : _GEN_7145; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7151 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_2 : _GEN_4781; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7152 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_2 : _GEN_7151; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7153 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_2 : _GEN_7152; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7154 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_2 : _GEN_7153; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7159 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_3 : _GEN_4789; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7160 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_3 : _GEN_7159; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7161 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_3 : _GEN_7160; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7162 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_3 : _GEN_7161; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7167 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_4 : _GEN_4797; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7168 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_4 : _GEN_7167; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7169 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_4 : _GEN_7168; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7170 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_4 : _GEN_7169; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7175 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_5 : _GEN_4805; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7176 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_5 : _GEN_7175; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7177 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_5 : _GEN_7176; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7178 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_5 : _GEN_7177; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7183 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_6 : _GEN_4813; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7184 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_6 : _GEN_7183; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7185 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_6 : _GEN_7184; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7186 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_6 : _GEN_7185; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7191 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_1_7 : _GEN_4821; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7192 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_2_7 : _GEN_7191; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7193 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_3_7 : _GEN_7192; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7194 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_5_4_7 : _GEN_7193; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7199 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_0 : _GEN_4829; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7200 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_0 : _GEN_7199; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7201 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_0 : _GEN_7200; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7202 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_0 : _GEN_7201; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7207 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_1 : _GEN_4837; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7208 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_1 : _GEN_7207; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7209 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_1 : _GEN_7208; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7210 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_1 : _GEN_7209; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7215 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_2 : _GEN_4845; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7216 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_2 : _GEN_7215; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7217 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_2 : _GEN_7216; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7218 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_2 : _GEN_7217; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7223 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_3 : _GEN_4853; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7224 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_3 : _GEN_7223; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7225 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_3 : _GEN_7224; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7226 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_3 : _GEN_7225; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7231 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_4 : _GEN_4861; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7232 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_4 : _GEN_7231; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7233 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_4 : _GEN_7232; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7234 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_4 : _GEN_7233; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7239 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_5 : _GEN_4869; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7240 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_5 : _GEN_7239; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7241 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_5 : _GEN_7240; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7242 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_5 : _GEN_7241; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7247 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_6 : _GEN_4877; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7248 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_6 : _GEN_7247; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7249 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_6 : _GEN_7248; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7250 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_6 : _GEN_7249; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7255 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_1_7 : _GEN_4885; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7256 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_2_7 : _GEN_7255; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7257 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_3_7 : _GEN_7256; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7258 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_6_4_7 : _GEN_7257; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7263 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_0 : _GEN_4893; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7264 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_0 : _GEN_7263; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7265 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_0 : _GEN_7264; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7266 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_0 : _GEN_7265; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7271 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_1 : _GEN_4901; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7272 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_1 : _GEN_7271; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7273 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_1 : _GEN_7272; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7274 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_1 : _GEN_7273; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7279 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_2 : _GEN_4909; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7280 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_2 : _GEN_7279; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7281 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_2 : _GEN_7280; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7282 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_2 : _GEN_7281; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7287 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_3 : _GEN_4917; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7288 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_3 : _GEN_7287; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7289 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_3 : _GEN_7288; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7290 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_3 : _GEN_7289; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7295 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_4 : _GEN_4925; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7296 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_4 : _GEN_7295; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7297 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_4 : _GEN_7296; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7298 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_4 : _GEN_7297; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7303 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_5 : _GEN_4933; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7304 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_5 : _GEN_7303; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7305 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_5 : _GEN_7304; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7306 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_5 : _GEN_7305; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7311 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_6 : _GEN_4941; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7312 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_6 : _GEN_7311; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7313 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_6 : _GEN_7312; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7314 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_6 : _GEN_7313; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7319 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_1_7 : _GEN_4949; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7320 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_2_7 : _GEN_7319; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7321 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_3_7 : _GEN_7320; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7322 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_7_4_7 : _GEN_7321; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7327 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_0 : _GEN_4957; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7328 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_0 : _GEN_7327; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7329 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_0 : _GEN_7328; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7330 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_0 : _GEN_7329; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7335 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_1 : _GEN_4965; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7336 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_1 : _GEN_7335; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7337 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_1 : _GEN_7336; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7338 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_1 : _GEN_7337; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7343 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_2 : _GEN_4973; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7344 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_2 : _GEN_7343; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7345 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_2 : _GEN_7344; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7346 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_2 : _GEN_7345; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7351 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_3 : _GEN_4981; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7352 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_3 : _GEN_7351; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7353 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_3 : _GEN_7352; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7354 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_3 : _GEN_7353; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7359 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_4 : _GEN_4989; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7360 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_4 : _GEN_7359; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7361 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_4 : _GEN_7360; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7362 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_4 : _GEN_7361; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7367 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_5 : _GEN_4997; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7368 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_5 : _GEN_7367; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7369 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_5 : _GEN_7368; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7370 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_5 : _GEN_7369; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7375 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_6 : _GEN_5005; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7376 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_6 : _GEN_7375; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7377 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_6 : _GEN_7376; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7378 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_6 : _GEN_7377; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7383 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_1_7 : _GEN_5013; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7384 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_2_7 : _GEN_7383; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7385 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_3_7 : _GEN_7384; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7386 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_8_4_7 : _GEN_7385; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7391 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_0 : _GEN_5021; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7392 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_0 : _GEN_7391; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7393 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_0 : _GEN_7392; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7394 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_0 : _GEN_7393; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7399 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_1 : _GEN_5029; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7400 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_1 : _GEN_7399; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7401 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_1 : _GEN_7400; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7402 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_1 : _GEN_7401; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7407 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_2 : _GEN_5037; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7408 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_2 : _GEN_7407; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7409 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_2 : _GEN_7408; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7410 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_2 : _GEN_7409; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7415 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_3 : _GEN_5045; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7416 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_3 : _GEN_7415; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7417 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_3 : _GEN_7416; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7418 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_3 : _GEN_7417; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7423 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_4 : _GEN_5053; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7424 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_4 : _GEN_7423; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7425 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_4 : _GEN_7424; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7426 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_4 : _GEN_7425; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7431 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_5 : _GEN_5061; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7432 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_5 : _GEN_7431; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7433 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_5 : _GEN_7432; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7434 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_5 : _GEN_7433; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7439 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_6 : _GEN_5069; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7440 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_6 : _GEN_7439; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7441 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_6 : _GEN_7440; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7442 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_6 : _GEN_7441; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7447 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_1_7 : _GEN_5077; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7448 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_2_7 : _GEN_7447; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7449 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_3_7 : _GEN_7448; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7450 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_9_4_7 : _GEN_7449; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7455 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_0 : _GEN_5085; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7456 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_0 : _GEN_7455; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7457 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_0 : _GEN_7456; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7458 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_0 : _GEN_7457; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7463 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_1 : _GEN_5093; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7464 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_1 : _GEN_7463; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7465 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_1 : _GEN_7464; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7466 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_1 : _GEN_7465; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7471 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_2 : _GEN_5101; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7472 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_2 : _GEN_7471; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7473 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_2 : _GEN_7472; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7474 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_2 : _GEN_7473; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7479 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_3 : _GEN_5109; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7480 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_3 : _GEN_7479; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7481 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_3 : _GEN_7480; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7482 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_3 : _GEN_7481; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7487 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_4 : _GEN_5117; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7488 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_4 : _GEN_7487; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7489 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_4 : _GEN_7488; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7490 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_4 : _GEN_7489; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7495 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_5 : _GEN_5125; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7496 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_5 : _GEN_7495; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7497 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_5 : _GEN_7496; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7498 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_5 : _GEN_7497; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7503 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_6 : _GEN_5133; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7504 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_6 : _GEN_7503; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7505 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_6 : _GEN_7504; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7506 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_6 : _GEN_7505; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7511 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_1_7 : _GEN_5141; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7512 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_2_7 : _GEN_7511; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7513 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_3_7 : _GEN_7512; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7514 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_10_4_7 : _GEN_7513; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7519 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_0 : _GEN_5149; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7520 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_0 : _GEN_7519; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7521 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_0 : _GEN_7520; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7522 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_0 : _GEN_7521; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7527 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_1 : _GEN_5157; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7528 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_1 : _GEN_7527; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7529 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_1 : _GEN_7528; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7530 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_1 : _GEN_7529; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7535 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_2 : _GEN_5165; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7536 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_2 : _GEN_7535; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7537 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_2 : _GEN_7536; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7538 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_2 : _GEN_7537; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7543 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_3 : _GEN_5173; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7544 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_3 : _GEN_7543; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7545 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_3 : _GEN_7544; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7546 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_3 : _GEN_7545; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7551 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_4 : _GEN_5181; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7552 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_4 : _GEN_7551; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7553 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_4 : _GEN_7552; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7554 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_4 : _GEN_7553; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7559 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_5 : _GEN_5189; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7560 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_5 : _GEN_7559; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7561 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_5 : _GEN_7560; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7562 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_5 : _GEN_7561; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7567 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_6 : _GEN_5197; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7568 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_6 : _GEN_7567; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7569 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_6 : _GEN_7568; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7570 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_6 : _GEN_7569; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7575 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_1_7 : _GEN_5205; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7576 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_2_7 : _GEN_7575; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7577 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_3_7 : _GEN_7576; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7578 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_11_4_7 : _GEN_7577; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7583 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_0 : _GEN_5213; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7584 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_0 : _GEN_7583; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7585 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_0 : _GEN_7584; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7586 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_0 : _GEN_7585; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7591 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_1 : _GEN_5221; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7592 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_1 : _GEN_7591; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7593 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_1 : _GEN_7592; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7594 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_1 : _GEN_7593; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7599 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_2 : _GEN_5229; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7600 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_2 : _GEN_7599; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7601 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_2 : _GEN_7600; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7602 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_2 : _GEN_7601; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7607 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_3 : _GEN_5237; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7608 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_3 : _GEN_7607; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7609 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_3 : _GEN_7608; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7610 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_3 : _GEN_7609; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7615 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_4 : _GEN_5245; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7616 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_4 : _GEN_7615; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7617 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_4 : _GEN_7616; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7618 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_4 : _GEN_7617; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7623 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_5 : _GEN_5253; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7624 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_5 : _GEN_7623; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7625 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_5 : _GEN_7624; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7626 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_5 : _GEN_7625; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7631 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_6 : _GEN_5261; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7632 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_6 : _GEN_7631; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7633 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_6 : _GEN_7632; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7634 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_6 : _GEN_7633; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7639 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_1_7 : _GEN_5269; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7640 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_2_7 : _GEN_7639; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7641 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_3_7 : _GEN_7640; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7642 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_12_4_7 : _GEN_7641; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7647 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_0 : _GEN_5277; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7648 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_0 : _GEN_7647; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7649 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_0 : _GEN_7648; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7650 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_0 : _GEN_7649; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7655 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_1 : _GEN_5285; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7656 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_1 : _GEN_7655; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7657 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_1 : _GEN_7656; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7658 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_1 : _GEN_7657; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7663 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_2 : _GEN_5293; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7664 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_2 : _GEN_7663; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7665 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_2 : _GEN_7664; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7666 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_2 : _GEN_7665; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7671 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_3 : _GEN_5301; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7672 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_3 : _GEN_7671; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7673 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_3 : _GEN_7672; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7674 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_3 : _GEN_7673; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7679 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_4 : _GEN_5309; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7680 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_4 : _GEN_7679; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7681 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_4 : _GEN_7680; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7682 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_4 : _GEN_7681; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7687 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_5 : _GEN_5317; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7688 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_5 : _GEN_7687; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7689 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_5 : _GEN_7688; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7690 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_5 : _GEN_7689; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7695 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_6 : _GEN_5325; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7696 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_6 : _GEN_7695; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7697 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_6 : _GEN_7696; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7698 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_6 : _GEN_7697; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7703 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_1_7 : _GEN_5333; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7704 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_2_7 : _GEN_7703; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7705 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_3_7 : _GEN_7704; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7706 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_13_4_7 : _GEN_7705; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7711 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_0 : _GEN_5341; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7712 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_0 : _GEN_7711; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7713 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_0 : _GEN_7712; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7714 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_0 : _GEN_7713; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7719 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_1 : _GEN_5349; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7720 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_1 : _GEN_7719; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7721 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_1 : _GEN_7720; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7722 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_1 : _GEN_7721; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7727 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_2 : _GEN_5357; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7728 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_2 : _GEN_7727; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7729 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_2 : _GEN_7728; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7730 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_2 : _GEN_7729; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7735 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_3 : _GEN_5365; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7736 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_3 : _GEN_7735; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7737 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_3 : _GEN_7736; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7738 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_3 : _GEN_7737; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7743 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_4 : _GEN_5373; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7744 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_4 : _GEN_7743; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7745 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_4 : _GEN_7744; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7746 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_4 : _GEN_7745; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7751 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_5 : _GEN_5381; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7752 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_5 : _GEN_7751; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7753 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_5 : _GEN_7752; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7754 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_5 : _GEN_7753; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7759 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_6 : _GEN_5389; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7760 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_6 : _GEN_7759; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7761 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_6 : _GEN_7760; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7762 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_6 : _GEN_7761; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7767 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_1_7 : _GEN_5397; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7768 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_2_7 : _GEN_7767; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7769 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_3_7 : _GEN_7768; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7770 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_14_4_7 : _GEN_7769; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7775 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_0 : _GEN_5405; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7776 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_0 : _GEN_7775; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7777 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_0 : _GEN_7776; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7778 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_0 : _GEN_7777; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7783 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_1 : _GEN_5413; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7784 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_1 : _GEN_7783; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7785 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_1 : _GEN_7784; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7786 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_1 : _GEN_7785; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7791 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_2 : _GEN_5421; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7792 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_2 : _GEN_7791; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7793 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_2 : _GEN_7792; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7794 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_2 : _GEN_7793; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7799 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_3 : _GEN_5429; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7800 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_3 : _GEN_7799; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7801 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_3 : _GEN_7800; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7802 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_3 : _GEN_7801; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7807 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_4 : _GEN_5437; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7808 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_4 : _GEN_7807; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7809 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_4 : _GEN_7808; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7810 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_4 : _GEN_7809; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7815 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_5 : _GEN_5445; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7816 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_5 : _GEN_7815; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7817 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_5 : _GEN_7816; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7818 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_5 : _GEN_7817; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7823 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_6 : _GEN_5453; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7824 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_6 : _GEN_7823; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7825 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_6 : _GEN_7824; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7826 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_6 : _GEN_7825; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7831 = 3'h1 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_1_7 : _GEN_5461; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7832 = 3'h2 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_2_7 : _GEN_7831; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7833 = 3'h3 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_3_7 : _GEN_7832; // @[Sbuffer.scala 824:{14,14}]
  wire [7:0] _GEN_7834 = 3'h4 == io_forward_1_paddr[5:3] ? dataModule_io_dataOut_15_4_7 : _GEN_7833; // @[Sbuffer.scala 824:{14,14}]
  reg [7:0] forward_data_candidate_reg_1_0_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_0_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_1_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_2_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_3_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_4_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_5_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_6_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_7_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_8_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_9_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_10_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_11_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_12_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_13_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_14_7; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_0; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_1; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_2; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_3; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_4; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_5; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_6; // @[Reg.scala 19:16]
  reg [7:0] forward_data_candidate_reg_1_15_7; // @[Reg.scala 19:16]
  wire  _selectedValidMask_T_263 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_0; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_0 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_0 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_0 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_0 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_0 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_0 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_0 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_0 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_0 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_0 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_0 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_0 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_0 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_0 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_0 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_0 |
    _selectedValidMask_T_263; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_294 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_1; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_1 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_1 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_1 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_1 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_1 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_1 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_1 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_1 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_1 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_1 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_1 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_1 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_1 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_1 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_1 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_1 |
    _selectedValidMask_T_294; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_325 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_2; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_2 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_2 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_2 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_2 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_2 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_2 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_2 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_2 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_2 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_2 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_2 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_2 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_2 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_2 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_2 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_2 |
    _selectedValidMask_T_325; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_356 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_3; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_3 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_3 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_3 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_3 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_3 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_3 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_3 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_3 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_3 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_3 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_3 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_3 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_3 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_3 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_3 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_3 |
    _selectedValidMask_T_356; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_387 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_4; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_4 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_4 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_4 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_4 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_4 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_4 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_4 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_4 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_4 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_4 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_4 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_4 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_4 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_4 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_4 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_4 |
    _selectedValidMask_T_387; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_418 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_5; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_5 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_5 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_5 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_5 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_5 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_5 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_5 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_5 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_5 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_5 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_5 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_5 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_5 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_5 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_5 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_5 |
    _selectedValidMask_T_418; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_449 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_6; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_6 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_6 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_6 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_6 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_6 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_6 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_6 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_6 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_6 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_6 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_6 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_6 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_6 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_6 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_6 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_6 |
    _selectedValidMask_T_449; // @[Mux.scala 27:73]
  wire  _selectedValidMask_T_480 = valid_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_7; // @[Mux.scala 27:73]
  wire  selectedValidMask_1_7 = valid_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_7 | valid_tag_match_reg_1_1 &
    forward_mask_candidate_reg_1_1_7 | valid_tag_match_reg_2_1 & forward_mask_candidate_reg_1_2_7 |
    valid_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_7 | valid_tag_match_reg_4_1 &
    forward_mask_candidate_reg_1_4_7 | valid_tag_match_reg_5_1 & forward_mask_candidate_reg_1_5_7 |
    valid_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_7 | valid_tag_match_reg_7_1 &
    forward_mask_candidate_reg_1_7_7 | valid_tag_match_reg_8_1 & forward_mask_candidate_reg_1_8_7 |
    valid_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_7 | valid_tag_match_reg_10_1 &
    forward_mask_candidate_reg_1_10_7 | valid_tag_match_reg_11_1 & forward_mask_candidate_reg_1_11_7 |
    valid_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_7 | valid_tag_match_reg_13_1 &
    forward_mask_candidate_reg_1_13_7 | valid_tag_match_reg_14_1 & forward_mask_candidate_reg_1_14_7 |
    _selectedValidMask_T_480; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_248 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_249 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_250 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_251 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_252 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_253 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_254 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_255 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_256 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_257 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_258 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_259 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_260 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_261 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_262 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_263 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_264 = _selectedValidData_T_248 | _selectedValidData_T_249; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_265 = _selectedValidData_T_264 | _selectedValidData_T_250; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_266 = _selectedValidData_T_265 | _selectedValidData_T_251; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_267 = _selectedValidData_T_266 | _selectedValidData_T_252; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_268 = _selectedValidData_T_267 | _selectedValidData_T_253; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_269 = _selectedValidData_T_268 | _selectedValidData_T_254; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_270 = _selectedValidData_T_269 | _selectedValidData_T_255; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_271 = _selectedValidData_T_270 | _selectedValidData_T_256; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_272 = _selectedValidData_T_271 | _selectedValidData_T_257; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_273 = _selectedValidData_T_272 | _selectedValidData_T_258; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_274 = _selectedValidData_T_273 | _selectedValidData_T_259; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_275 = _selectedValidData_T_274 | _selectedValidData_T_260; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_276 = _selectedValidData_T_275 | _selectedValidData_T_261; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_277 = _selectedValidData_T_276 | _selectedValidData_T_262; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_0 = _selectedValidData_T_277 | _selectedValidData_T_263; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_279 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_280 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_281 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_282 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_283 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_284 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_285 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_286 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_287 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_288 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_289 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_290 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_291 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_292 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_293 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_294 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_295 = _selectedValidData_T_279 | _selectedValidData_T_280; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_296 = _selectedValidData_T_295 | _selectedValidData_T_281; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_297 = _selectedValidData_T_296 | _selectedValidData_T_282; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_298 = _selectedValidData_T_297 | _selectedValidData_T_283; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_299 = _selectedValidData_T_298 | _selectedValidData_T_284; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_300 = _selectedValidData_T_299 | _selectedValidData_T_285; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_301 = _selectedValidData_T_300 | _selectedValidData_T_286; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_302 = _selectedValidData_T_301 | _selectedValidData_T_287; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_303 = _selectedValidData_T_302 | _selectedValidData_T_288; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_304 = _selectedValidData_T_303 | _selectedValidData_T_289; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_305 = _selectedValidData_T_304 | _selectedValidData_T_290; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_306 = _selectedValidData_T_305 | _selectedValidData_T_291; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_307 = _selectedValidData_T_306 | _selectedValidData_T_292; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_308 = _selectedValidData_T_307 | _selectedValidData_T_293; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_1 = _selectedValidData_T_308 | _selectedValidData_T_294; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_310 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_311 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_312 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_313 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_314 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_315 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_316 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_317 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_318 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_319 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_320 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_321 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_322 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_323 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_324 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_325 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_326 = _selectedValidData_T_310 | _selectedValidData_T_311; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_327 = _selectedValidData_T_326 | _selectedValidData_T_312; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_328 = _selectedValidData_T_327 | _selectedValidData_T_313; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_329 = _selectedValidData_T_328 | _selectedValidData_T_314; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_330 = _selectedValidData_T_329 | _selectedValidData_T_315; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_331 = _selectedValidData_T_330 | _selectedValidData_T_316; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_332 = _selectedValidData_T_331 | _selectedValidData_T_317; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_333 = _selectedValidData_T_332 | _selectedValidData_T_318; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_334 = _selectedValidData_T_333 | _selectedValidData_T_319; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_335 = _selectedValidData_T_334 | _selectedValidData_T_320; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_336 = _selectedValidData_T_335 | _selectedValidData_T_321; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_337 = _selectedValidData_T_336 | _selectedValidData_T_322; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_338 = _selectedValidData_T_337 | _selectedValidData_T_323; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_339 = _selectedValidData_T_338 | _selectedValidData_T_324; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_2 = _selectedValidData_T_339 | _selectedValidData_T_325; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_341 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_342 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_343 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_344 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_345 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_346 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_347 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_348 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_349 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_350 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_351 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_352 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_353 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_354 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_355 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_356 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_357 = _selectedValidData_T_341 | _selectedValidData_T_342; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_358 = _selectedValidData_T_357 | _selectedValidData_T_343; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_359 = _selectedValidData_T_358 | _selectedValidData_T_344; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_360 = _selectedValidData_T_359 | _selectedValidData_T_345; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_361 = _selectedValidData_T_360 | _selectedValidData_T_346; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_362 = _selectedValidData_T_361 | _selectedValidData_T_347; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_363 = _selectedValidData_T_362 | _selectedValidData_T_348; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_364 = _selectedValidData_T_363 | _selectedValidData_T_349; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_365 = _selectedValidData_T_364 | _selectedValidData_T_350; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_366 = _selectedValidData_T_365 | _selectedValidData_T_351; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_367 = _selectedValidData_T_366 | _selectedValidData_T_352; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_368 = _selectedValidData_T_367 | _selectedValidData_T_353; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_369 = _selectedValidData_T_368 | _selectedValidData_T_354; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_370 = _selectedValidData_T_369 | _selectedValidData_T_355; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_3 = _selectedValidData_T_370 | _selectedValidData_T_356; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_372 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_373 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_374 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_375 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_376 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_377 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_378 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_379 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_380 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_381 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_382 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_383 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_384 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_385 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_386 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_387 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_388 = _selectedValidData_T_372 | _selectedValidData_T_373; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_389 = _selectedValidData_T_388 | _selectedValidData_T_374; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_390 = _selectedValidData_T_389 | _selectedValidData_T_375; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_391 = _selectedValidData_T_390 | _selectedValidData_T_376; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_392 = _selectedValidData_T_391 | _selectedValidData_T_377; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_393 = _selectedValidData_T_392 | _selectedValidData_T_378; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_394 = _selectedValidData_T_393 | _selectedValidData_T_379; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_395 = _selectedValidData_T_394 | _selectedValidData_T_380; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_396 = _selectedValidData_T_395 | _selectedValidData_T_381; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_397 = _selectedValidData_T_396 | _selectedValidData_T_382; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_398 = _selectedValidData_T_397 | _selectedValidData_T_383; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_399 = _selectedValidData_T_398 | _selectedValidData_T_384; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_400 = _selectedValidData_T_399 | _selectedValidData_T_385; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_401 = _selectedValidData_T_400 | _selectedValidData_T_386; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_4 = _selectedValidData_T_401 | _selectedValidData_T_387; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_403 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_404 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_405 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_406 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_407 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_408 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_409 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_410 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_411 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_412 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_413 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_414 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_415 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_416 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_417 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_418 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_419 = _selectedValidData_T_403 | _selectedValidData_T_404; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_420 = _selectedValidData_T_419 | _selectedValidData_T_405; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_421 = _selectedValidData_T_420 | _selectedValidData_T_406; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_422 = _selectedValidData_T_421 | _selectedValidData_T_407; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_423 = _selectedValidData_T_422 | _selectedValidData_T_408; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_424 = _selectedValidData_T_423 | _selectedValidData_T_409; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_425 = _selectedValidData_T_424 | _selectedValidData_T_410; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_426 = _selectedValidData_T_425 | _selectedValidData_T_411; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_427 = _selectedValidData_T_426 | _selectedValidData_T_412; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_428 = _selectedValidData_T_427 | _selectedValidData_T_413; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_429 = _selectedValidData_T_428 | _selectedValidData_T_414; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_430 = _selectedValidData_T_429 | _selectedValidData_T_415; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_431 = _selectedValidData_T_430 | _selectedValidData_T_416; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_432 = _selectedValidData_T_431 | _selectedValidData_T_417; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_5 = _selectedValidData_T_432 | _selectedValidData_T_418; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_434 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_435 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_436 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_437 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_438 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_439 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_440 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_441 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_442 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_443 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_444 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_445 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_446 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_447 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_448 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_449 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_450 = _selectedValidData_T_434 | _selectedValidData_T_435; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_451 = _selectedValidData_T_450 | _selectedValidData_T_436; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_452 = _selectedValidData_T_451 | _selectedValidData_T_437; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_453 = _selectedValidData_T_452 | _selectedValidData_T_438; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_454 = _selectedValidData_T_453 | _selectedValidData_T_439; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_455 = _selectedValidData_T_454 | _selectedValidData_T_440; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_456 = _selectedValidData_T_455 | _selectedValidData_T_441; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_457 = _selectedValidData_T_456 | _selectedValidData_T_442; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_458 = _selectedValidData_T_457 | _selectedValidData_T_443; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_459 = _selectedValidData_T_458 | _selectedValidData_T_444; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_460 = _selectedValidData_T_459 | _selectedValidData_T_445; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_461 = _selectedValidData_T_460 | _selectedValidData_T_446; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_462 = _selectedValidData_T_461 | _selectedValidData_T_447; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_463 = _selectedValidData_T_462 | _selectedValidData_T_448; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_6 = _selectedValidData_T_463 | _selectedValidData_T_449; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_465 = valid_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_466 = valid_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_467 = valid_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_468 = valid_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_469 = valid_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_470 = valid_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_471 = valid_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_472 = valid_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_473 = valid_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_474 = valid_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_475 = valid_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_476 = valid_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_477 = valid_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_478 = valid_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_479 = valid_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_480 = valid_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_481 = _selectedValidData_T_465 | _selectedValidData_T_466; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_482 = _selectedValidData_T_481 | _selectedValidData_T_467; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_483 = _selectedValidData_T_482 | _selectedValidData_T_468; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_484 = _selectedValidData_T_483 | _selectedValidData_T_469; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_485 = _selectedValidData_T_484 | _selectedValidData_T_470; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_486 = _selectedValidData_T_485 | _selectedValidData_T_471; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_487 = _selectedValidData_T_486 | _selectedValidData_T_472; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_488 = _selectedValidData_T_487 | _selectedValidData_T_473; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_489 = _selectedValidData_T_488 | _selectedValidData_T_474; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_490 = _selectedValidData_T_489 | _selectedValidData_T_475; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_491 = _selectedValidData_T_490 | _selectedValidData_T_476; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_492 = _selectedValidData_T_491 | _selectedValidData_T_477; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_493 = _selectedValidData_T_492 | _selectedValidData_T_478; // @[Mux.scala 27:73]
  wire [7:0] _selectedValidData_T_494 = _selectedValidData_T_493 | _selectedValidData_T_479; // @[Mux.scala 27:73]
  wire [7:0] selectedValidData_1_7 = _selectedValidData_T_494 | _selectedValidData_T_480; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_263 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_0; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_0 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_0 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_0 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_0 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_0 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_0 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_0 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_0 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_0 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_0 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_0 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_0 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_0 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_0 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_0 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_0 | _selectedInflightMask_T_263; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_294 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_1; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_1 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_1 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_1 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_1 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_1 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_1 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_1 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_1 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_1 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_1 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_1 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_1 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_1 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_1 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_1 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_1 | _selectedInflightMask_T_294; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_325 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_2; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_2 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_2 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_2 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_2 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_2 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_2 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_2 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_2 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_2 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_2 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_2 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_2 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_2 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_2 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_2 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_2 | _selectedInflightMask_T_325; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_356 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_3; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_3 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_3 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_3 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_3 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_3 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_3 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_3 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_3 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_3 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_3 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_3 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_3 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_3 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_3 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_3 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_3 | _selectedInflightMask_T_356; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_387 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_4; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_4 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_4 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_4 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_4 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_4 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_4 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_4 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_4 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_4 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_4 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_4 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_4 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_4 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_4 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_4 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_4 | _selectedInflightMask_T_387; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_418 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_5; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_5 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_5 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_5 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_5 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_5 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_5 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_5 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_5 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_5 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_5 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_5 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_5 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_5 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_5 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_5 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_5 | _selectedInflightMask_T_418; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_449 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_6; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_6 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_6 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_6 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_6 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_6 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_6 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_6 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_6 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_6 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_6 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_6 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_6 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_6 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_6 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_6 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_6 | _selectedInflightMask_T_449; // @[Mux.scala 27:73]
  wire  _selectedInflightMask_T_480 = inflight_tag_match_reg_15_1 & forward_mask_candidate_reg_1_15_7; // @[Mux.scala 27:73]
  wire  selectedInflightMask_1_7 = inflight_tag_match_reg_0_1 & forward_mask_candidate_reg_1_0_7 |
    inflight_tag_match_reg_1_1 & forward_mask_candidate_reg_1_1_7 | inflight_tag_match_reg_2_1 &
    forward_mask_candidate_reg_1_2_7 | inflight_tag_match_reg_3_1 & forward_mask_candidate_reg_1_3_7 |
    inflight_tag_match_reg_4_1 & forward_mask_candidate_reg_1_4_7 | inflight_tag_match_reg_5_1 &
    forward_mask_candidate_reg_1_5_7 | inflight_tag_match_reg_6_1 & forward_mask_candidate_reg_1_6_7 |
    inflight_tag_match_reg_7_1 & forward_mask_candidate_reg_1_7_7 | inflight_tag_match_reg_8_1 &
    forward_mask_candidate_reg_1_8_7 | inflight_tag_match_reg_9_1 & forward_mask_candidate_reg_1_9_7 |
    inflight_tag_match_reg_10_1 & forward_mask_candidate_reg_1_10_7 | inflight_tag_match_reg_11_1 &
    forward_mask_candidate_reg_1_11_7 | inflight_tag_match_reg_12_1 & forward_mask_candidate_reg_1_12_7 |
    inflight_tag_match_reg_13_1 & forward_mask_candidate_reg_1_13_7 | inflight_tag_match_reg_14_1 &
    forward_mask_candidate_reg_1_14_7 | _selectedInflightMask_T_480; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_248 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_249 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_250 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_251 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_252 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_253 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_254 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_255 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_256 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_257 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_258 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_259 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_260 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_261 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_262 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_263 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_264 = _selectedInflightData_T_248 | _selectedInflightData_T_249; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_265 = _selectedInflightData_T_264 | _selectedInflightData_T_250; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_266 = _selectedInflightData_T_265 | _selectedInflightData_T_251; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_267 = _selectedInflightData_T_266 | _selectedInflightData_T_252; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_268 = _selectedInflightData_T_267 | _selectedInflightData_T_253; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_269 = _selectedInflightData_T_268 | _selectedInflightData_T_254; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_270 = _selectedInflightData_T_269 | _selectedInflightData_T_255; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_271 = _selectedInflightData_T_270 | _selectedInflightData_T_256; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_272 = _selectedInflightData_T_271 | _selectedInflightData_T_257; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_273 = _selectedInflightData_T_272 | _selectedInflightData_T_258; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_274 = _selectedInflightData_T_273 | _selectedInflightData_T_259; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_275 = _selectedInflightData_T_274 | _selectedInflightData_T_260; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_276 = _selectedInflightData_T_275 | _selectedInflightData_T_261; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_277 = _selectedInflightData_T_276 | _selectedInflightData_T_262; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_0 = _selectedInflightData_T_277 | _selectedInflightData_T_263; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_279 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_280 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_281 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_282 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_283 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_284 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_285 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_286 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_287 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_288 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_289 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_290 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_291 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_292 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_293 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_294 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_295 = _selectedInflightData_T_279 | _selectedInflightData_T_280; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_296 = _selectedInflightData_T_295 | _selectedInflightData_T_281; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_297 = _selectedInflightData_T_296 | _selectedInflightData_T_282; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_298 = _selectedInflightData_T_297 | _selectedInflightData_T_283; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_299 = _selectedInflightData_T_298 | _selectedInflightData_T_284; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_300 = _selectedInflightData_T_299 | _selectedInflightData_T_285; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_301 = _selectedInflightData_T_300 | _selectedInflightData_T_286; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_302 = _selectedInflightData_T_301 | _selectedInflightData_T_287; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_303 = _selectedInflightData_T_302 | _selectedInflightData_T_288; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_304 = _selectedInflightData_T_303 | _selectedInflightData_T_289; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_305 = _selectedInflightData_T_304 | _selectedInflightData_T_290; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_306 = _selectedInflightData_T_305 | _selectedInflightData_T_291; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_307 = _selectedInflightData_T_306 | _selectedInflightData_T_292; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_308 = _selectedInflightData_T_307 | _selectedInflightData_T_293; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_1 = _selectedInflightData_T_308 | _selectedInflightData_T_294; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_310 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_311 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_312 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_313 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_314 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_315 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_316 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_317 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_318 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_319 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_320 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_321 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_322 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_323 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_324 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_325 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_326 = _selectedInflightData_T_310 | _selectedInflightData_T_311; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_327 = _selectedInflightData_T_326 | _selectedInflightData_T_312; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_328 = _selectedInflightData_T_327 | _selectedInflightData_T_313; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_329 = _selectedInflightData_T_328 | _selectedInflightData_T_314; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_330 = _selectedInflightData_T_329 | _selectedInflightData_T_315; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_331 = _selectedInflightData_T_330 | _selectedInflightData_T_316; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_332 = _selectedInflightData_T_331 | _selectedInflightData_T_317; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_333 = _selectedInflightData_T_332 | _selectedInflightData_T_318; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_334 = _selectedInflightData_T_333 | _selectedInflightData_T_319; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_335 = _selectedInflightData_T_334 | _selectedInflightData_T_320; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_336 = _selectedInflightData_T_335 | _selectedInflightData_T_321; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_337 = _selectedInflightData_T_336 | _selectedInflightData_T_322; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_338 = _selectedInflightData_T_337 | _selectedInflightData_T_323; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_339 = _selectedInflightData_T_338 | _selectedInflightData_T_324; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_2 = _selectedInflightData_T_339 | _selectedInflightData_T_325; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_341 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_342 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_343 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_344 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_345 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_346 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_347 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_348 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_349 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_350 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_351 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_352 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_353 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_354 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_355 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_356 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_3 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_357 = _selectedInflightData_T_341 | _selectedInflightData_T_342; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_358 = _selectedInflightData_T_357 | _selectedInflightData_T_343; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_359 = _selectedInflightData_T_358 | _selectedInflightData_T_344; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_360 = _selectedInflightData_T_359 | _selectedInflightData_T_345; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_361 = _selectedInflightData_T_360 | _selectedInflightData_T_346; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_362 = _selectedInflightData_T_361 | _selectedInflightData_T_347; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_363 = _selectedInflightData_T_362 | _selectedInflightData_T_348; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_364 = _selectedInflightData_T_363 | _selectedInflightData_T_349; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_365 = _selectedInflightData_T_364 | _selectedInflightData_T_350; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_366 = _selectedInflightData_T_365 | _selectedInflightData_T_351; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_367 = _selectedInflightData_T_366 | _selectedInflightData_T_352; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_368 = _selectedInflightData_T_367 | _selectedInflightData_T_353; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_369 = _selectedInflightData_T_368 | _selectedInflightData_T_354; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_370 = _selectedInflightData_T_369 | _selectedInflightData_T_355; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_3 = _selectedInflightData_T_370 | _selectedInflightData_T_356; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_372 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_373 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_374 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_375 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_376 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_377 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_378 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_379 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_380 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_381 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_382 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_383 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_384 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_385 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_386 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_387 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_4 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_388 = _selectedInflightData_T_372 | _selectedInflightData_T_373; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_389 = _selectedInflightData_T_388 | _selectedInflightData_T_374; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_390 = _selectedInflightData_T_389 | _selectedInflightData_T_375; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_391 = _selectedInflightData_T_390 | _selectedInflightData_T_376; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_392 = _selectedInflightData_T_391 | _selectedInflightData_T_377; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_393 = _selectedInflightData_T_392 | _selectedInflightData_T_378; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_394 = _selectedInflightData_T_393 | _selectedInflightData_T_379; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_395 = _selectedInflightData_T_394 | _selectedInflightData_T_380; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_396 = _selectedInflightData_T_395 | _selectedInflightData_T_381; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_397 = _selectedInflightData_T_396 | _selectedInflightData_T_382; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_398 = _selectedInflightData_T_397 | _selectedInflightData_T_383; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_399 = _selectedInflightData_T_398 | _selectedInflightData_T_384; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_400 = _selectedInflightData_T_399 | _selectedInflightData_T_385; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_401 = _selectedInflightData_T_400 | _selectedInflightData_T_386; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_4 = _selectedInflightData_T_401 | _selectedInflightData_T_387; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_403 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_404 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_405 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_406 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_407 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_408 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_409 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_410 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_411 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_412 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_413 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_414 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_415 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_416 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_417 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_418 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_5 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_419 = _selectedInflightData_T_403 | _selectedInflightData_T_404; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_420 = _selectedInflightData_T_419 | _selectedInflightData_T_405; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_421 = _selectedInflightData_T_420 | _selectedInflightData_T_406; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_422 = _selectedInflightData_T_421 | _selectedInflightData_T_407; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_423 = _selectedInflightData_T_422 | _selectedInflightData_T_408; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_424 = _selectedInflightData_T_423 | _selectedInflightData_T_409; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_425 = _selectedInflightData_T_424 | _selectedInflightData_T_410; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_426 = _selectedInflightData_T_425 | _selectedInflightData_T_411; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_427 = _selectedInflightData_T_426 | _selectedInflightData_T_412; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_428 = _selectedInflightData_T_427 | _selectedInflightData_T_413; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_429 = _selectedInflightData_T_428 | _selectedInflightData_T_414; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_430 = _selectedInflightData_T_429 | _selectedInflightData_T_415; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_431 = _selectedInflightData_T_430 | _selectedInflightData_T_416; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_432 = _selectedInflightData_T_431 | _selectedInflightData_T_417; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_5 = _selectedInflightData_T_432 | _selectedInflightData_T_418; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_434 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_435 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_436 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_437 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_438 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_439 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_440 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_441 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_442 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_443 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_444 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_445 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_446 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_447 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_448 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_449 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_6 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_450 = _selectedInflightData_T_434 | _selectedInflightData_T_435; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_451 = _selectedInflightData_T_450 | _selectedInflightData_T_436; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_452 = _selectedInflightData_T_451 | _selectedInflightData_T_437; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_453 = _selectedInflightData_T_452 | _selectedInflightData_T_438; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_454 = _selectedInflightData_T_453 | _selectedInflightData_T_439; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_455 = _selectedInflightData_T_454 | _selectedInflightData_T_440; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_456 = _selectedInflightData_T_455 | _selectedInflightData_T_441; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_457 = _selectedInflightData_T_456 | _selectedInflightData_T_442; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_458 = _selectedInflightData_T_457 | _selectedInflightData_T_443; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_459 = _selectedInflightData_T_458 | _selectedInflightData_T_444; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_460 = _selectedInflightData_T_459 | _selectedInflightData_T_445; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_461 = _selectedInflightData_T_460 | _selectedInflightData_T_446; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_462 = _selectedInflightData_T_461 | _selectedInflightData_T_447; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_463 = _selectedInflightData_T_462 | _selectedInflightData_T_448; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_6 = _selectedInflightData_T_463 | _selectedInflightData_T_449; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_465 = inflight_tag_match_reg_0_1 ? forward_data_candidate_reg_1_0_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_466 = inflight_tag_match_reg_1_1 ? forward_data_candidate_reg_1_1_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_467 = inflight_tag_match_reg_2_1 ? forward_data_candidate_reg_1_2_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_468 = inflight_tag_match_reg_3_1 ? forward_data_candidate_reg_1_3_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_469 = inflight_tag_match_reg_4_1 ? forward_data_candidate_reg_1_4_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_470 = inflight_tag_match_reg_5_1 ? forward_data_candidate_reg_1_5_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_471 = inflight_tag_match_reg_6_1 ? forward_data_candidate_reg_1_6_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_472 = inflight_tag_match_reg_7_1 ? forward_data_candidate_reg_1_7_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_473 = inflight_tag_match_reg_8_1 ? forward_data_candidate_reg_1_8_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_474 = inflight_tag_match_reg_9_1 ? forward_data_candidate_reg_1_9_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_475 = inflight_tag_match_reg_10_1 ? forward_data_candidate_reg_1_10_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_476 = inflight_tag_match_reg_11_1 ? forward_data_candidate_reg_1_11_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_477 = inflight_tag_match_reg_12_1 ? forward_data_candidate_reg_1_12_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_478 = inflight_tag_match_reg_13_1 ? forward_data_candidate_reg_1_13_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_479 = inflight_tag_match_reg_14_1 ? forward_data_candidate_reg_1_14_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_480 = inflight_tag_match_reg_15_1 ? forward_data_candidate_reg_1_15_7 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_481 = _selectedInflightData_T_465 | _selectedInflightData_T_466; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_482 = _selectedInflightData_T_481 | _selectedInflightData_T_467; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_483 = _selectedInflightData_T_482 | _selectedInflightData_T_468; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_484 = _selectedInflightData_T_483 | _selectedInflightData_T_469; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_485 = _selectedInflightData_T_484 | _selectedInflightData_T_470; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_486 = _selectedInflightData_T_485 | _selectedInflightData_T_471; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_487 = _selectedInflightData_T_486 | _selectedInflightData_T_472; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_488 = _selectedInflightData_T_487 | _selectedInflightData_T_473; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_489 = _selectedInflightData_T_488 | _selectedInflightData_T_474; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_490 = _selectedInflightData_T_489 | _selectedInflightData_T_475; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_491 = _selectedInflightData_T_490 | _selectedInflightData_T_476; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_492 = _selectedInflightData_T_491 | _selectedInflightData_T_477; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_493 = _selectedInflightData_T_492 | _selectedInflightData_T_478; // @[Mux.scala 27:73]
  wire [7:0] _selectedInflightData_T_494 = _selectedInflightData_T_493 | _selectedInflightData_T_479; // @[Mux.scala 27:73]
  wire [7:0] selectedInflightData_1_7 = _selectedInflightData_T_494 | _selectedInflightData_T_480; // @[Mux.scala 27:73]
  wire  _perf_valid_entry_count_T_1 = ~invalidMask_0; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_3 = ~invalidMask_1; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_5 = ~invalidMask_2; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_7 = ~invalidMask_3; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_9 = ~invalidMask_4; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_11 = ~invalidMask_5; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_13 = ~invalidMask_6; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_15 = ~invalidMask_7; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_17 = ~invalidMask_8; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_19 = ~invalidMask_9; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_21 = ~invalidMask_10; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_23 = ~invalidMask_11; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_25 = ~invalidMask_12; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_27 = ~invalidMask_13; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_29 = ~invalidMask_14; // @[Sbuffer.scala 873:75]
  wire  _perf_valid_entry_count_T_31 = ~invalidMask_15; // @[Sbuffer.scala 873:75]
  wire [7:0] perf_valid_entry_count_lo = {_perf_valid_entry_count_T_15,_perf_valid_entry_count_T_13,
    _perf_valid_entry_count_T_11,_perf_valid_entry_count_T_9,_perf_valid_entry_count_T_7,_perf_valid_entry_count_T_5,
    _perf_valid_entry_count_T_3,_perf_valid_entry_count_T_1}; // @[Sbuffer.scala 873:92]
  wire [15:0] _perf_valid_entry_count_T_32 = {_perf_valid_entry_count_T_31,_perf_valid_entry_count_T_29,
    _perf_valid_entry_count_T_27,_perf_valid_entry_count_T_25,_perf_valid_entry_count_T_23,_perf_valid_entry_count_T_21,
    _perf_valid_entry_count_T_19,_perf_valid_entry_count_T_17,perf_valid_entry_count_lo}; // @[Sbuffer.scala 873:92]
  wire [1:0] _perf_valid_entry_count_T_49 = _perf_valid_entry_count_T_32[0] + _perf_valid_entry_count_T_32[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_51 = _perf_valid_entry_count_T_32[2] + _perf_valid_entry_count_T_32[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _perf_valid_entry_count_T_53 = _perf_valid_entry_count_T_49 + _perf_valid_entry_count_T_51; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_55 = _perf_valid_entry_count_T_32[4] + _perf_valid_entry_count_T_32[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_57 = _perf_valid_entry_count_T_32[6] + _perf_valid_entry_count_T_32[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _perf_valid_entry_count_T_59 = _perf_valid_entry_count_T_55 + _perf_valid_entry_count_T_57; // @[Bitwise.scala 51:90]
  wire [3:0] _perf_valid_entry_count_T_61 = _perf_valid_entry_count_T_53 + _perf_valid_entry_count_T_59; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_63 = _perf_valid_entry_count_T_32[8] + _perf_valid_entry_count_T_32[9]; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_65 = _perf_valid_entry_count_T_32[10] + _perf_valid_entry_count_T_32[11]; // @[Bitwise.scala 51:90]
  wire [2:0] _perf_valid_entry_count_T_67 = _perf_valid_entry_count_T_63 + _perf_valid_entry_count_T_65; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_69 = _perf_valid_entry_count_T_32[12] + _perf_valid_entry_count_T_32[13]; // @[Bitwise.scala 51:90]
  wire [1:0] _perf_valid_entry_count_T_71 = _perf_valid_entry_count_T_32[14] + _perf_valid_entry_count_T_32[15]; // @[Bitwise.scala 51:90]
  wire [2:0] _perf_valid_entry_count_T_73 = _perf_valid_entry_count_T_69 + _perf_valid_entry_count_T_71; // @[Bitwise.scala 51:90]
  wire [3:0] _perf_valid_entry_count_T_75 = _perf_valid_entry_count_T_67 + _perf_valid_entry_count_T_73; // @[Bitwise.scala 51:90]
  reg [4:0] perf_valid_entry_count; // @[Sbuffer.scala 873:39]
  wire [1:0] _T_1099 = {io_in_1_valid,io_in_0_valid}; // @[Sbuffer.scala 896:65]
  wire [1:0] _T_1106 = {_dataModule_io_writeReq_1_valid_T,_dataModule_io_writeReq_0_valid_T}; // @[Sbuffer.scala 897:66]
  wire  _T_1112 = _dataModule_io_writeReq_0_valid_T & canMerge_0; // @[Sbuffer.scala 898:95]
  wire  _T_1114 = _dataModule_io_writeReq_1_valid_T & canMerge_1; // @[Sbuffer.scala 898:95]
  wire [1:0] _T_1115 = {_T_1114,_T_1112}; // @[Sbuffer.scala 898:113]
  wire  _T_1122 = _dataModule_io_writeReq_0_valid_T & ~canMerge_0; // @[Sbuffer.scala 899:95]
  wire  _T_1125 = _dataModule_io_writeReq_1_valid_T & ~canMerge_1; // @[Sbuffer.scala 899:95]
  wire [1:0] _T_1126 = {_T_1125,_T_1122}; // @[Sbuffer.scala 899:114]
  wire [4:0] _T_1135 = 5'h10 / 3'h4; // @[Sbuffer.scala 909:72]
  wire [4:0] _T_1139 = 5'h10 / 2'h2; // @[Sbuffer.scala 910:126]
  wire [6:0] _T_1144 = 5'h10 * 2'h3; // @[Sbuffer.scala 911:126]
  wire [6:0] _T_1145 = _T_1144 / 3'h4; // @[Sbuffer.scala 911:130]
  wire [6:0] _GEN_3180 = {{2'd0}, perf_valid_entry_count}; // @[Sbuffer.scala 911:105]
  reg [1:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg [1:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg [1:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg [1:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg [1:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg [1:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg [1:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg [1:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_4_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_5_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_6_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_7_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_8_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_8_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_9_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_9_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_10_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_10_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_11_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_11_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_12_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_12_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_13_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_13_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_14_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_14_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_15_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_15_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  reg  io_perf_16_value_REG; // @[PerfCounterUtils.scala 172:35]
  reg  io_perf_16_value_REG_1; // @[PerfCounterUtils.scala 172:27]
  SbufferData dataModule ( // @[Sbuffer.scala 270:26]
    .clock(dataModule_clock),
    .reset(dataModule_reset),
    .io_writeReq_0_valid(dataModule_io_writeReq_0_valid),
    .io_writeReq_0_bits_wvec(dataModule_io_writeReq_0_bits_wvec),
    .io_writeReq_0_bits_mask(dataModule_io_writeReq_0_bits_mask),
    .io_writeReq_0_bits_data(dataModule_io_writeReq_0_bits_data),
    .io_writeReq_0_bits_wordOffset(dataModule_io_writeReq_0_bits_wordOffset),
    .io_writeReq_0_bits_wline(dataModule_io_writeReq_0_bits_wline),
    .io_writeReq_1_valid(dataModule_io_writeReq_1_valid),
    .io_writeReq_1_bits_wvec(dataModule_io_writeReq_1_bits_wvec),
    .io_writeReq_1_bits_mask(dataModule_io_writeReq_1_bits_mask),
    .io_writeReq_1_bits_data(dataModule_io_writeReq_1_bits_data),
    .io_writeReq_1_bits_wordOffset(dataModule_io_writeReq_1_bits_wordOffset),
    .io_writeReq_1_bits_wline(dataModule_io_writeReq_1_bits_wline),
    .io_maskFlushReq_0_valid(dataModule_io_maskFlushReq_0_valid),
    .io_maskFlushReq_0_bits_wvec(dataModule_io_maskFlushReq_0_bits_wvec),
    .io_maskFlushReq_1_valid(dataModule_io_maskFlushReq_1_valid),
    .io_maskFlushReq_1_bits_wvec(dataModule_io_maskFlushReq_1_bits_wvec),
    .io_dataOut_0_0_0(dataModule_io_dataOut_0_0_0),
    .io_dataOut_0_0_1(dataModule_io_dataOut_0_0_1),
    .io_dataOut_0_0_2(dataModule_io_dataOut_0_0_2),
    .io_dataOut_0_0_3(dataModule_io_dataOut_0_0_3),
    .io_dataOut_0_0_4(dataModule_io_dataOut_0_0_4),
    .io_dataOut_0_0_5(dataModule_io_dataOut_0_0_5),
    .io_dataOut_0_0_6(dataModule_io_dataOut_0_0_6),
    .io_dataOut_0_0_7(dataModule_io_dataOut_0_0_7),
    .io_dataOut_0_1_0(dataModule_io_dataOut_0_1_0),
    .io_dataOut_0_1_1(dataModule_io_dataOut_0_1_1),
    .io_dataOut_0_1_2(dataModule_io_dataOut_0_1_2),
    .io_dataOut_0_1_3(dataModule_io_dataOut_0_1_3),
    .io_dataOut_0_1_4(dataModule_io_dataOut_0_1_4),
    .io_dataOut_0_1_5(dataModule_io_dataOut_0_1_5),
    .io_dataOut_0_1_6(dataModule_io_dataOut_0_1_6),
    .io_dataOut_0_1_7(dataModule_io_dataOut_0_1_7),
    .io_dataOut_0_2_0(dataModule_io_dataOut_0_2_0),
    .io_dataOut_0_2_1(dataModule_io_dataOut_0_2_1),
    .io_dataOut_0_2_2(dataModule_io_dataOut_0_2_2),
    .io_dataOut_0_2_3(dataModule_io_dataOut_0_2_3),
    .io_dataOut_0_2_4(dataModule_io_dataOut_0_2_4),
    .io_dataOut_0_2_5(dataModule_io_dataOut_0_2_5),
    .io_dataOut_0_2_6(dataModule_io_dataOut_0_2_6),
    .io_dataOut_0_2_7(dataModule_io_dataOut_0_2_7),
    .io_dataOut_0_3_0(dataModule_io_dataOut_0_3_0),
    .io_dataOut_0_3_1(dataModule_io_dataOut_0_3_1),
    .io_dataOut_0_3_2(dataModule_io_dataOut_0_3_2),
    .io_dataOut_0_3_3(dataModule_io_dataOut_0_3_3),
    .io_dataOut_0_3_4(dataModule_io_dataOut_0_3_4),
    .io_dataOut_0_3_5(dataModule_io_dataOut_0_3_5),
    .io_dataOut_0_3_6(dataModule_io_dataOut_0_3_6),
    .io_dataOut_0_3_7(dataModule_io_dataOut_0_3_7),
    .io_dataOut_0_4_0(dataModule_io_dataOut_0_4_0),
    .io_dataOut_0_4_1(dataModule_io_dataOut_0_4_1),
    .io_dataOut_0_4_2(dataModule_io_dataOut_0_4_2),
    .io_dataOut_0_4_3(dataModule_io_dataOut_0_4_3),
    .io_dataOut_0_4_4(dataModule_io_dataOut_0_4_4),
    .io_dataOut_0_4_5(dataModule_io_dataOut_0_4_5),
    .io_dataOut_0_4_6(dataModule_io_dataOut_0_4_6),
    .io_dataOut_0_4_7(dataModule_io_dataOut_0_4_7),
    .io_dataOut_0_5_0(dataModule_io_dataOut_0_5_0),
    .io_dataOut_0_5_1(dataModule_io_dataOut_0_5_1),
    .io_dataOut_0_5_2(dataModule_io_dataOut_0_5_2),
    .io_dataOut_0_5_3(dataModule_io_dataOut_0_5_3),
    .io_dataOut_0_5_4(dataModule_io_dataOut_0_5_4),
    .io_dataOut_0_5_5(dataModule_io_dataOut_0_5_5),
    .io_dataOut_0_5_6(dataModule_io_dataOut_0_5_6),
    .io_dataOut_0_5_7(dataModule_io_dataOut_0_5_7),
    .io_dataOut_0_6_0(dataModule_io_dataOut_0_6_0),
    .io_dataOut_0_6_1(dataModule_io_dataOut_0_6_1),
    .io_dataOut_0_6_2(dataModule_io_dataOut_0_6_2),
    .io_dataOut_0_6_3(dataModule_io_dataOut_0_6_3),
    .io_dataOut_0_6_4(dataModule_io_dataOut_0_6_4),
    .io_dataOut_0_6_5(dataModule_io_dataOut_0_6_5),
    .io_dataOut_0_6_6(dataModule_io_dataOut_0_6_6),
    .io_dataOut_0_6_7(dataModule_io_dataOut_0_6_7),
    .io_dataOut_0_7_0(dataModule_io_dataOut_0_7_0),
    .io_dataOut_0_7_1(dataModule_io_dataOut_0_7_1),
    .io_dataOut_0_7_2(dataModule_io_dataOut_0_7_2),
    .io_dataOut_0_7_3(dataModule_io_dataOut_0_7_3),
    .io_dataOut_0_7_4(dataModule_io_dataOut_0_7_4),
    .io_dataOut_0_7_5(dataModule_io_dataOut_0_7_5),
    .io_dataOut_0_7_6(dataModule_io_dataOut_0_7_6),
    .io_dataOut_0_7_7(dataModule_io_dataOut_0_7_7),
    .io_dataOut_1_0_0(dataModule_io_dataOut_1_0_0),
    .io_dataOut_1_0_1(dataModule_io_dataOut_1_0_1),
    .io_dataOut_1_0_2(dataModule_io_dataOut_1_0_2),
    .io_dataOut_1_0_3(dataModule_io_dataOut_1_0_3),
    .io_dataOut_1_0_4(dataModule_io_dataOut_1_0_4),
    .io_dataOut_1_0_5(dataModule_io_dataOut_1_0_5),
    .io_dataOut_1_0_6(dataModule_io_dataOut_1_0_6),
    .io_dataOut_1_0_7(dataModule_io_dataOut_1_0_7),
    .io_dataOut_1_1_0(dataModule_io_dataOut_1_1_0),
    .io_dataOut_1_1_1(dataModule_io_dataOut_1_1_1),
    .io_dataOut_1_1_2(dataModule_io_dataOut_1_1_2),
    .io_dataOut_1_1_3(dataModule_io_dataOut_1_1_3),
    .io_dataOut_1_1_4(dataModule_io_dataOut_1_1_4),
    .io_dataOut_1_1_5(dataModule_io_dataOut_1_1_5),
    .io_dataOut_1_1_6(dataModule_io_dataOut_1_1_6),
    .io_dataOut_1_1_7(dataModule_io_dataOut_1_1_7),
    .io_dataOut_1_2_0(dataModule_io_dataOut_1_2_0),
    .io_dataOut_1_2_1(dataModule_io_dataOut_1_2_1),
    .io_dataOut_1_2_2(dataModule_io_dataOut_1_2_2),
    .io_dataOut_1_2_3(dataModule_io_dataOut_1_2_3),
    .io_dataOut_1_2_4(dataModule_io_dataOut_1_2_4),
    .io_dataOut_1_2_5(dataModule_io_dataOut_1_2_5),
    .io_dataOut_1_2_6(dataModule_io_dataOut_1_2_6),
    .io_dataOut_1_2_7(dataModule_io_dataOut_1_2_7),
    .io_dataOut_1_3_0(dataModule_io_dataOut_1_3_0),
    .io_dataOut_1_3_1(dataModule_io_dataOut_1_3_1),
    .io_dataOut_1_3_2(dataModule_io_dataOut_1_3_2),
    .io_dataOut_1_3_3(dataModule_io_dataOut_1_3_3),
    .io_dataOut_1_3_4(dataModule_io_dataOut_1_3_4),
    .io_dataOut_1_3_5(dataModule_io_dataOut_1_3_5),
    .io_dataOut_1_3_6(dataModule_io_dataOut_1_3_6),
    .io_dataOut_1_3_7(dataModule_io_dataOut_1_3_7),
    .io_dataOut_1_4_0(dataModule_io_dataOut_1_4_0),
    .io_dataOut_1_4_1(dataModule_io_dataOut_1_4_1),
    .io_dataOut_1_4_2(dataModule_io_dataOut_1_4_2),
    .io_dataOut_1_4_3(dataModule_io_dataOut_1_4_3),
    .io_dataOut_1_4_4(dataModule_io_dataOut_1_4_4),
    .io_dataOut_1_4_5(dataModule_io_dataOut_1_4_5),
    .io_dataOut_1_4_6(dataModule_io_dataOut_1_4_6),
    .io_dataOut_1_4_7(dataModule_io_dataOut_1_4_7),
    .io_dataOut_1_5_0(dataModule_io_dataOut_1_5_0),
    .io_dataOut_1_5_1(dataModule_io_dataOut_1_5_1),
    .io_dataOut_1_5_2(dataModule_io_dataOut_1_5_2),
    .io_dataOut_1_5_3(dataModule_io_dataOut_1_5_3),
    .io_dataOut_1_5_4(dataModule_io_dataOut_1_5_4),
    .io_dataOut_1_5_5(dataModule_io_dataOut_1_5_5),
    .io_dataOut_1_5_6(dataModule_io_dataOut_1_5_6),
    .io_dataOut_1_5_7(dataModule_io_dataOut_1_5_7),
    .io_dataOut_1_6_0(dataModule_io_dataOut_1_6_0),
    .io_dataOut_1_6_1(dataModule_io_dataOut_1_6_1),
    .io_dataOut_1_6_2(dataModule_io_dataOut_1_6_2),
    .io_dataOut_1_6_3(dataModule_io_dataOut_1_6_3),
    .io_dataOut_1_6_4(dataModule_io_dataOut_1_6_4),
    .io_dataOut_1_6_5(dataModule_io_dataOut_1_6_5),
    .io_dataOut_1_6_6(dataModule_io_dataOut_1_6_6),
    .io_dataOut_1_6_7(dataModule_io_dataOut_1_6_7),
    .io_dataOut_1_7_0(dataModule_io_dataOut_1_7_0),
    .io_dataOut_1_7_1(dataModule_io_dataOut_1_7_1),
    .io_dataOut_1_7_2(dataModule_io_dataOut_1_7_2),
    .io_dataOut_1_7_3(dataModule_io_dataOut_1_7_3),
    .io_dataOut_1_7_4(dataModule_io_dataOut_1_7_4),
    .io_dataOut_1_7_5(dataModule_io_dataOut_1_7_5),
    .io_dataOut_1_7_6(dataModule_io_dataOut_1_7_6),
    .io_dataOut_1_7_7(dataModule_io_dataOut_1_7_7),
    .io_dataOut_2_0_0(dataModule_io_dataOut_2_0_0),
    .io_dataOut_2_0_1(dataModule_io_dataOut_2_0_1),
    .io_dataOut_2_0_2(dataModule_io_dataOut_2_0_2),
    .io_dataOut_2_0_3(dataModule_io_dataOut_2_0_3),
    .io_dataOut_2_0_4(dataModule_io_dataOut_2_0_4),
    .io_dataOut_2_0_5(dataModule_io_dataOut_2_0_5),
    .io_dataOut_2_0_6(dataModule_io_dataOut_2_0_6),
    .io_dataOut_2_0_7(dataModule_io_dataOut_2_0_7),
    .io_dataOut_2_1_0(dataModule_io_dataOut_2_1_0),
    .io_dataOut_2_1_1(dataModule_io_dataOut_2_1_1),
    .io_dataOut_2_1_2(dataModule_io_dataOut_2_1_2),
    .io_dataOut_2_1_3(dataModule_io_dataOut_2_1_3),
    .io_dataOut_2_1_4(dataModule_io_dataOut_2_1_4),
    .io_dataOut_2_1_5(dataModule_io_dataOut_2_1_5),
    .io_dataOut_2_1_6(dataModule_io_dataOut_2_1_6),
    .io_dataOut_2_1_7(dataModule_io_dataOut_2_1_7),
    .io_dataOut_2_2_0(dataModule_io_dataOut_2_2_0),
    .io_dataOut_2_2_1(dataModule_io_dataOut_2_2_1),
    .io_dataOut_2_2_2(dataModule_io_dataOut_2_2_2),
    .io_dataOut_2_2_3(dataModule_io_dataOut_2_2_3),
    .io_dataOut_2_2_4(dataModule_io_dataOut_2_2_4),
    .io_dataOut_2_2_5(dataModule_io_dataOut_2_2_5),
    .io_dataOut_2_2_6(dataModule_io_dataOut_2_2_6),
    .io_dataOut_2_2_7(dataModule_io_dataOut_2_2_7),
    .io_dataOut_2_3_0(dataModule_io_dataOut_2_3_0),
    .io_dataOut_2_3_1(dataModule_io_dataOut_2_3_1),
    .io_dataOut_2_3_2(dataModule_io_dataOut_2_3_2),
    .io_dataOut_2_3_3(dataModule_io_dataOut_2_3_3),
    .io_dataOut_2_3_4(dataModule_io_dataOut_2_3_4),
    .io_dataOut_2_3_5(dataModule_io_dataOut_2_3_5),
    .io_dataOut_2_3_6(dataModule_io_dataOut_2_3_6),
    .io_dataOut_2_3_7(dataModule_io_dataOut_2_3_7),
    .io_dataOut_2_4_0(dataModule_io_dataOut_2_4_0),
    .io_dataOut_2_4_1(dataModule_io_dataOut_2_4_1),
    .io_dataOut_2_4_2(dataModule_io_dataOut_2_4_2),
    .io_dataOut_2_4_3(dataModule_io_dataOut_2_4_3),
    .io_dataOut_2_4_4(dataModule_io_dataOut_2_4_4),
    .io_dataOut_2_4_5(dataModule_io_dataOut_2_4_5),
    .io_dataOut_2_4_6(dataModule_io_dataOut_2_4_6),
    .io_dataOut_2_4_7(dataModule_io_dataOut_2_4_7),
    .io_dataOut_2_5_0(dataModule_io_dataOut_2_5_0),
    .io_dataOut_2_5_1(dataModule_io_dataOut_2_5_1),
    .io_dataOut_2_5_2(dataModule_io_dataOut_2_5_2),
    .io_dataOut_2_5_3(dataModule_io_dataOut_2_5_3),
    .io_dataOut_2_5_4(dataModule_io_dataOut_2_5_4),
    .io_dataOut_2_5_5(dataModule_io_dataOut_2_5_5),
    .io_dataOut_2_5_6(dataModule_io_dataOut_2_5_6),
    .io_dataOut_2_5_7(dataModule_io_dataOut_2_5_7),
    .io_dataOut_2_6_0(dataModule_io_dataOut_2_6_0),
    .io_dataOut_2_6_1(dataModule_io_dataOut_2_6_1),
    .io_dataOut_2_6_2(dataModule_io_dataOut_2_6_2),
    .io_dataOut_2_6_3(dataModule_io_dataOut_2_6_3),
    .io_dataOut_2_6_4(dataModule_io_dataOut_2_6_4),
    .io_dataOut_2_6_5(dataModule_io_dataOut_2_6_5),
    .io_dataOut_2_6_6(dataModule_io_dataOut_2_6_6),
    .io_dataOut_2_6_7(dataModule_io_dataOut_2_6_7),
    .io_dataOut_2_7_0(dataModule_io_dataOut_2_7_0),
    .io_dataOut_2_7_1(dataModule_io_dataOut_2_7_1),
    .io_dataOut_2_7_2(dataModule_io_dataOut_2_7_2),
    .io_dataOut_2_7_3(dataModule_io_dataOut_2_7_3),
    .io_dataOut_2_7_4(dataModule_io_dataOut_2_7_4),
    .io_dataOut_2_7_5(dataModule_io_dataOut_2_7_5),
    .io_dataOut_2_7_6(dataModule_io_dataOut_2_7_6),
    .io_dataOut_2_7_7(dataModule_io_dataOut_2_7_7),
    .io_dataOut_3_0_0(dataModule_io_dataOut_3_0_0),
    .io_dataOut_3_0_1(dataModule_io_dataOut_3_0_1),
    .io_dataOut_3_0_2(dataModule_io_dataOut_3_0_2),
    .io_dataOut_3_0_3(dataModule_io_dataOut_3_0_3),
    .io_dataOut_3_0_4(dataModule_io_dataOut_3_0_4),
    .io_dataOut_3_0_5(dataModule_io_dataOut_3_0_5),
    .io_dataOut_3_0_6(dataModule_io_dataOut_3_0_6),
    .io_dataOut_3_0_7(dataModule_io_dataOut_3_0_7),
    .io_dataOut_3_1_0(dataModule_io_dataOut_3_1_0),
    .io_dataOut_3_1_1(dataModule_io_dataOut_3_1_1),
    .io_dataOut_3_1_2(dataModule_io_dataOut_3_1_2),
    .io_dataOut_3_1_3(dataModule_io_dataOut_3_1_3),
    .io_dataOut_3_1_4(dataModule_io_dataOut_3_1_4),
    .io_dataOut_3_1_5(dataModule_io_dataOut_3_1_5),
    .io_dataOut_3_1_6(dataModule_io_dataOut_3_1_6),
    .io_dataOut_3_1_7(dataModule_io_dataOut_3_1_7),
    .io_dataOut_3_2_0(dataModule_io_dataOut_3_2_0),
    .io_dataOut_3_2_1(dataModule_io_dataOut_3_2_1),
    .io_dataOut_3_2_2(dataModule_io_dataOut_3_2_2),
    .io_dataOut_3_2_3(dataModule_io_dataOut_3_2_3),
    .io_dataOut_3_2_4(dataModule_io_dataOut_3_2_4),
    .io_dataOut_3_2_5(dataModule_io_dataOut_3_2_5),
    .io_dataOut_3_2_6(dataModule_io_dataOut_3_2_6),
    .io_dataOut_3_2_7(dataModule_io_dataOut_3_2_7),
    .io_dataOut_3_3_0(dataModule_io_dataOut_3_3_0),
    .io_dataOut_3_3_1(dataModule_io_dataOut_3_3_1),
    .io_dataOut_3_3_2(dataModule_io_dataOut_3_3_2),
    .io_dataOut_3_3_3(dataModule_io_dataOut_3_3_3),
    .io_dataOut_3_3_4(dataModule_io_dataOut_3_3_4),
    .io_dataOut_3_3_5(dataModule_io_dataOut_3_3_5),
    .io_dataOut_3_3_6(dataModule_io_dataOut_3_3_6),
    .io_dataOut_3_3_7(dataModule_io_dataOut_3_3_7),
    .io_dataOut_3_4_0(dataModule_io_dataOut_3_4_0),
    .io_dataOut_3_4_1(dataModule_io_dataOut_3_4_1),
    .io_dataOut_3_4_2(dataModule_io_dataOut_3_4_2),
    .io_dataOut_3_4_3(dataModule_io_dataOut_3_4_3),
    .io_dataOut_3_4_4(dataModule_io_dataOut_3_4_4),
    .io_dataOut_3_4_5(dataModule_io_dataOut_3_4_5),
    .io_dataOut_3_4_6(dataModule_io_dataOut_3_4_6),
    .io_dataOut_3_4_7(dataModule_io_dataOut_3_4_7),
    .io_dataOut_3_5_0(dataModule_io_dataOut_3_5_0),
    .io_dataOut_3_5_1(dataModule_io_dataOut_3_5_1),
    .io_dataOut_3_5_2(dataModule_io_dataOut_3_5_2),
    .io_dataOut_3_5_3(dataModule_io_dataOut_3_5_3),
    .io_dataOut_3_5_4(dataModule_io_dataOut_3_5_4),
    .io_dataOut_3_5_5(dataModule_io_dataOut_3_5_5),
    .io_dataOut_3_5_6(dataModule_io_dataOut_3_5_6),
    .io_dataOut_3_5_7(dataModule_io_dataOut_3_5_7),
    .io_dataOut_3_6_0(dataModule_io_dataOut_3_6_0),
    .io_dataOut_3_6_1(dataModule_io_dataOut_3_6_1),
    .io_dataOut_3_6_2(dataModule_io_dataOut_3_6_2),
    .io_dataOut_3_6_3(dataModule_io_dataOut_3_6_3),
    .io_dataOut_3_6_4(dataModule_io_dataOut_3_6_4),
    .io_dataOut_3_6_5(dataModule_io_dataOut_3_6_5),
    .io_dataOut_3_6_6(dataModule_io_dataOut_3_6_6),
    .io_dataOut_3_6_7(dataModule_io_dataOut_3_6_7),
    .io_dataOut_3_7_0(dataModule_io_dataOut_3_7_0),
    .io_dataOut_3_7_1(dataModule_io_dataOut_3_7_1),
    .io_dataOut_3_7_2(dataModule_io_dataOut_3_7_2),
    .io_dataOut_3_7_3(dataModule_io_dataOut_3_7_3),
    .io_dataOut_3_7_4(dataModule_io_dataOut_3_7_4),
    .io_dataOut_3_7_5(dataModule_io_dataOut_3_7_5),
    .io_dataOut_3_7_6(dataModule_io_dataOut_3_7_6),
    .io_dataOut_3_7_7(dataModule_io_dataOut_3_7_7),
    .io_dataOut_4_0_0(dataModule_io_dataOut_4_0_0),
    .io_dataOut_4_0_1(dataModule_io_dataOut_4_0_1),
    .io_dataOut_4_0_2(dataModule_io_dataOut_4_0_2),
    .io_dataOut_4_0_3(dataModule_io_dataOut_4_0_3),
    .io_dataOut_4_0_4(dataModule_io_dataOut_4_0_4),
    .io_dataOut_4_0_5(dataModule_io_dataOut_4_0_5),
    .io_dataOut_4_0_6(dataModule_io_dataOut_4_0_6),
    .io_dataOut_4_0_7(dataModule_io_dataOut_4_0_7),
    .io_dataOut_4_1_0(dataModule_io_dataOut_4_1_0),
    .io_dataOut_4_1_1(dataModule_io_dataOut_4_1_1),
    .io_dataOut_4_1_2(dataModule_io_dataOut_4_1_2),
    .io_dataOut_4_1_3(dataModule_io_dataOut_4_1_3),
    .io_dataOut_4_1_4(dataModule_io_dataOut_4_1_4),
    .io_dataOut_4_1_5(dataModule_io_dataOut_4_1_5),
    .io_dataOut_4_1_6(dataModule_io_dataOut_4_1_6),
    .io_dataOut_4_1_7(dataModule_io_dataOut_4_1_7),
    .io_dataOut_4_2_0(dataModule_io_dataOut_4_2_0),
    .io_dataOut_4_2_1(dataModule_io_dataOut_4_2_1),
    .io_dataOut_4_2_2(dataModule_io_dataOut_4_2_2),
    .io_dataOut_4_2_3(dataModule_io_dataOut_4_2_3),
    .io_dataOut_4_2_4(dataModule_io_dataOut_4_2_4),
    .io_dataOut_4_2_5(dataModule_io_dataOut_4_2_5),
    .io_dataOut_4_2_6(dataModule_io_dataOut_4_2_6),
    .io_dataOut_4_2_7(dataModule_io_dataOut_4_2_7),
    .io_dataOut_4_3_0(dataModule_io_dataOut_4_3_0),
    .io_dataOut_4_3_1(dataModule_io_dataOut_4_3_1),
    .io_dataOut_4_3_2(dataModule_io_dataOut_4_3_2),
    .io_dataOut_4_3_3(dataModule_io_dataOut_4_3_3),
    .io_dataOut_4_3_4(dataModule_io_dataOut_4_3_4),
    .io_dataOut_4_3_5(dataModule_io_dataOut_4_3_5),
    .io_dataOut_4_3_6(dataModule_io_dataOut_4_3_6),
    .io_dataOut_4_3_7(dataModule_io_dataOut_4_3_7),
    .io_dataOut_4_4_0(dataModule_io_dataOut_4_4_0),
    .io_dataOut_4_4_1(dataModule_io_dataOut_4_4_1),
    .io_dataOut_4_4_2(dataModule_io_dataOut_4_4_2),
    .io_dataOut_4_4_3(dataModule_io_dataOut_4_4_3),
    .io_dataOut_4_4_4(dataModule_io_dataOut_4_4_4),
    .io_dataOut_4_4_5(dataModule_io_dataOut_4_4_5),
    .io_dataOut_4_4_6(dataModule_io_dataOut_4_4_6),
    .io_dataOut_4_4_7(dataModule_io_dataOut_4_4_7),
    .io_dataOut_4_5_0(dataModule_io_dataOut_4_5_0),
    .io_dataOut_4_5_1(dataModule_io_dataOut_4_5_1),
    .io_dataOut_4_5_2(dataModule_io_dataOut_4_5_2),
    .io_dataOut_4_5_3(dataModule_io_dataOut_4_5_3),
    .io_dataOut_4_5_4(dataModule_io_dataOut_4_5_4),
    .io_dataOut_4_5_5(dataModule_io_dataOut_4_5_5),
    .io_dataOut_4_5_6(dataModule_io_dataOut_4_5_6),
    .io_dataOut_4_5_7(dataModule_io_dataOut_4_5_7),
    .io_dataOut_4_6_0(dataModule_io_dataOut_4_6_0),
    .io_dataOut_4_6_1(dataModule_io_dataOut_4_6_1),
    .io_dataOut_4_6_2(dataModule_io_dataOut_4_6_2),
    .io_dataOut_4_6_3(dataModule_io_dataOut_4_6_3),
    .io_dataOut_4_6_4(dataModule_io_dataOut_4_6_4),
    .io_dataOut_4_6_5(dataModule_io_dataOut_4_6_5),
    .io_dataOut_4_6_6(dataModule_io_dataOut_4_6_6),
    .io_dataOut_4_6_7(dataModule_io_dataOut_4_6_7),
    .io_dataOut_4_7_0(dataModule_io_dataOut_4_7_0),
    .io_dataOut_4_7_1(dataModule_io_dataOut_4_7_1),
    .io_dataOut_4_7_2(dataModule_io_dataOut_4_7_2),
    .io_dataOut_4_7_3(dataModule_io_dataOut_4_7_3),
    .io_dataOut_4_7_4(dataModule_io_dataOut_4_7_4),
    .io_dataOut_4_7_5(dataModule_io_dataOut_4_7_5),
    .io_dataOut_4_7_6(dataModule_io_dataOut_4_7_6),
    .io_dataOut_4_7_7(dataModule_io_dataOut_4_7_7),
    .io_dataOut_5_0_0(dataModule_io_dataOut_5_0_0),
    .io_dataOut_5_0_1(dataModule_io_dataOut_5_0_1),
    .io_dataOut_5_0_2(dataModule_io_dataOut_5_0_2),
    .io_dataOut_5_0_3(dataModule_io_dataOut_5_0_3),
    .io_dataOut_5_0_4(dataModule_io_dataOut_5_0_4),
    .io_dataOut_5_0_5(dataModule_io_dataOut_5_0_5),
    .io_dataOut_5_0_6(dataModule_io_dataOut_5_0_6),
    .io_dataOut_5_0_7(dataModule_io_dataOut_5_0_7),
    .io_dataOut_5_1_0(dataModule_io_dataOut_5_1_0),
    .io_dataOut_5_1_1(dataModule_io_dataOut_5_1_1),
    .io_dataOut_5_1_2(dataModule_io_dataOut_5_1_2),
    .io_dataOut_5_1_3(dataModule_io_dataOut_5_1_3),
    .io_dataOut_5_1_4(dataModule_io_dataOut_5_1_4),
    .io_dataOut_5_1_5(dataModule_io_dataOut_5_1_5),
    .io_dataOut_5_1_6(dataModule_io_dataOut_5_1_6),
    .io_dataOut_5_1_7(dataModule_io_dataOut_5_1_7),
    .io_dataOut_5_2_0(dataModule_io_dataOut_5_2_0),
    .io_dataOut_5_2_1(dataModule_io_dataOut_5_2_1),
    .io_dataOut_5_2_2(dataModule_io_dataOut_5_2_2),
    .io_dataOut_5_2_3(dataModule_io_dataOut_5_2_3),
    .io_dataOut_5_2_4(dataModule_io_dataOut_5_2_4),
    .io_dataOut_5_2_5(dataModule_io_dataOut_5_2_5),
    .io_dataOut_5_2_6(dataModule_io_dataOut_5_2_6),
    .io_dataOut_5_2_7(dataModule_io_dataOut_5_2_7),
    .io_dataOut_5_3_0(dataModule_io_dataOut_5_3_0),
    .io_dataOut_5_3_1(dataModule_io_dataOut_5_3_1),
    .io_dataOut_5_3_2(dataModule_io_dataOut_5_3_2),
    .io_dataOut_5_3_3(dataModule_io_dataOut_5_3_3),
    .io_dataOut_5_3_4(dataModule_io_dataOut_5_3_4),
    .io_dataOut_5_3_5(dataModule_io_dataOut_5_3_5),
    .io_dataOut_5_3_6(dataModule_io_dataOut_5_3_6),
    .io_dataOut_5_3_7(dataModule_io_dataOut_5_3_7),
    .io_dataOut_5_4_0(dataModule_io_dataOut_5_4_0),
    .io_dataOut_5_4_1(dataModule_io_dataOut_5_4_1),
    .io_dataOut_5_4_2(dataModule_io_dataOut_5_4_2),
    .io_dataOut_5_4_3(dataModule_io_dataOut_5_4_3),
    .io_dataOut_5_4_4(dataModule_io_dataOut_5_4_4),
    .io_dataOut_5_4_5(dataModule_io_dataOut_5_4_5),
    .io_dataOut_5_4_6(dataModule_io_dataOut_5_4_6),
    .io_dataOut_5_4_7(dataModule_io_dataOut_5_4_7),
    .io_dataOut_5_5_0(dataModule_io_dataOut_5_5_0),
    .io_dataOut_5_5_1(dataModule_io_dataOut_5_5_1),
    .io_dataOut_5_5_2(dataModule_io_dataOut_5_5_2),
    .io_dataOut_5_5_3(dataModule_io_dataOut_5_5_3),
    .io_dataOut_5_5_4(dataModule_io_dataOut_5_5_4),
    .io_dataOut_5_5_5(dataModule_io_dataOut_5_5_5),
    .io_dataOut_5_5_6(dataModule_io_dataOut_5_5_6),
    .io_dataOut_5_5_7(dataModule_io_dataOut_5_5_7),
    .io_dataOut_5_6_0(dataModule_io_dataOut_5_6_0),
    .io_dataOut_5_6_1(dataModule_io_dataOut_5_6_1),
    .io_dataOut_5_6_2(dataModule_io_dataOut_5_6_2),
    .io_dataOut_5_6_3(dataModule_io_dataOut_5_6_3),
    .io_dataOut_5_6_4(dataModule_io_dataOut_5_6_4),
    .io_dataOut_5_6_5(dataModule_io_dataOut_5_6_5),
    .io_dataOut_5_6_6(dataModule_io_dataOut_5_6_6),
    .io_dataOut_5_6_7(dataModule_io_dataOut_5_6_7),
    .io_dataOut_5_7_0(dataModule_io_dataOut_5_7_0),
    .io_dataOut_5_7_1(dataModule_io_dataOut_5_7_1),
    .io_dataOut_5_7_2(dataModule_io_dataOut_5_7_2),
    .io_dataOut_5_7_3(dataModule_io_dataOut_5_7_3),
    .io_dataOut_5_7_4(dataModule_io_dataOut_5_7_4),
    .io_dataOut_5_7_5(dataModule_io_dataOut_5_7_5),
    .io_dataOut_5_7_6(dataModule_io_dataOut_5_7_6),
    .io_dataOut_5_7_7(dataModule_io_dataOut_5_7_7),
    .io_dataOut_6_0_0(dataModule_io_dataOut_6_0_0),
    .io_dataOut_6_0_1(dataModule_io_dataOut_6_0_1),
    .io_dataOut_6_0_2(dataModule_io_dataOut_6_0_2),
    .io_dataOut_6_0_3(dataModule_io_dataOut_6_0_3),
    .io_dataOut_6_0_4(dataModule_io_dataOut_6_0_4),
    .io_dataOut_6_0_5(dataModule_io_dataOut_6_0_5),
    .io_dataOut_6_0_6(dataModule_io_dataOut_6_0_6),
    .io_dataOut_6_0_7(dataModule_io_dataOut_6_0_7),
    .io_dataOut_6_1_0(dataModule_io_dataOut_6_1_0),
    .io_dataOut_6_1_1(dataModule_io_dataOut_6_1_1),
    .io_dataOut_6_1_2(dataModule_io_dataOut_6_1_2),
    .io_dataOut_6_1_3(dataModule_io_dataOut_6_1_3),
    .io_dataOut_6_1_4(dataModule_io_dataOut_6_1_4),
    .io_dataOut_6_1_5(dataModule_io_dataOut_6_1_5),
    .io_dataOut_6_1_6(dataModule_io_dataOut_6_1_6),
    .io_dataOut_6_1_7(dataModule_io_dataOut_6_1_7),
    .io_dataOut_6_2_0(dataModule_io_dataOut_6_2_0),
    .io_dataOut_6_2_1(dataModule_io_dataOut_6_2_1),
    .io_dataOut_6_2_2(dataModule_io_dataOut_6_2_2),
    .io_dataOut_6_2_3(dataModule_io_dataOut_6_2_3),
    .io_dataOut_6_2_4(dataModule_io_dataOut_6_2_4),
    .io_dataOut_6_2_5(dataModule_io_dataOut_6_2_5),
    .io_dataOut_6_2_6(dataModule_io_dataOut_6_2_6),
    .io_dataOut_6_2_7(dataModule_io_dataOut_6_2_7),
    .io_dataOut_6_3_0(dataModule_io_dataOut_6_3_0),
    .io_dataOut_6_3_1(dataModule_io_dataOut_6_3_1),
    .io_dataOut_6_3_2(dataModule_io_dataOut_6_3_2),
    .io_dataOut_6_3_3(dataModule_io_dataOut_6_3_3),
    .io_dataOut_6_3_4(dataModule_io_dataOut_6_3_4),
    .io_dataOut_6_3_5(dataModule_io_dataOut_6_3_5),
    .io_dataOut_6_3_6(dataModule_io_dataOut_6_3_6),
    .io_dataOut_6_3_7(dataModule_io_dataOut_6_3_7),
    .io_dataOut_6_4_0(dataModule_io_dataOut_6_4_0),
    .io_dataOut_6_4_1(dataModule_io_dataOut_6_4_1),
    .io_dataOut_6_4_2(dataModule_io_dataOut_6_4_2),
    .io_dataOut_6_4_3(dataModule_io_dataOut_6_4_3),
    .io_dataOut_6_4_4(dataModule_io_dataOut_6_4_4),
    .io_dataOut_6_4_5(dataModule_io_dataOut_6_4_5),
    .io_dataOut_6_4_6(dataModule_io_dataOut_6_4_6),
    .io_dataOut_6_4_7(dataModule_io_dataOut_6_4_7),
    .io_dataOut_6_5_0(dataModule_io_dataOut_6_5_0),
    .io_dataOut_6_5_1(dataModule_io_dataOut_6_5_1),
    .io_dataOut_6_5_2(dataModule_io_dataOut_6_5_2),
    .io_dataOut_6_5_3(dataModule_io_dataOut_6_5_3),
    .io_dataOut_6_5_4(dataModule_io_dataOut_6_5_4),
    .io_dataOut_6_5_5(dataModule_io_dataOut_6_5_5),
    .io_dataOut_6_5_6(dataModule_io_dataOut_6_5_6),
    .io_dataOut_6_5_7(dataModule_io_dataOut_6_5_7),
    .io_dataOut_6_6_0(dataModule_io_dataOut_6_6_0),
    .io_dataOut_6_6_1(dataModule_io_dataOut_6_6_1),
    .io_dataOut_6_6_2(dataModule_io_dataOut_6_6_2),
    .io_dataOut_6_6_3(dataModule_io_dataOut_6_6_3),
    .io_dataOut_6_6_4(dataModule_io_dataOut_6_6_4),
    .io_dataOut_6_6_5(dataModule_io_dataOut_6_6_5),
    .io_dataOut_6_6_6(dataModule_io_dataOut_6_6_6),
    .io_dataOut_6_6_7(dataModule_io_dataOut_6_6_7),
    .io_dataOut_6_7_0(dataModule_io_dataOut_6_7_0),
    .io_dataOut_6_7_1(dataModule_io_dataOut_6_7_1),
    .io_dataOut_6_7_2(dataModule_io_dataOut_6_7_2),
    .io_dataOut_6_7_3(dataModule_io_dataOut_6_7_3),
    .io_dataOut_6_7_4(dataModule_io_dataOut_6_7_4),
    .io_dataOut_6_7_5(dataModule_io_dataOut_6_7_5),
    .io_dataOut_6_7_6(dataModule_io_dataOut_6_7_6),
    .io_dataOut_6_7_7(dataModule_io_dataOut_6_7_7),
    .io_dataOut_7_0_0(dataModule_io_dataOut_7_0_0),
    .io_dataOut_7_0_1(dataModule_io_dataOut_7_0_1),
    .io_dataOut_7_0_2(dataModule_io_dataOut_7_0_2),
    .io_dataOut_7_0_3(dataModule_io_dataOut_7_0_3),
    .io_dataOut_7_0_4(dataModule_io_dataOut_7_0_4),
    .io_dataOut_7_0_5(dataModule_io_dataOut_7_0_5),
    .io_dataOut_7_0_6(dataModule_io_dataOut_7_0_6),
    .io_dataOut_7_0_7(dataModule_io_dataOut_7_0_7),
    .io_dataOut_7_1_0(dataModule_io_dataOut_7_1_0),
    .io_dataOut_7_1_1(dataModule_io_dataOut_7_1_1),
    .io_dataOut_7_1_2(dataModule_io_dataOut_7_1_2),
    .io_dataOut_7_1_3(dataModule_io_dataOut_7_1_3),
    .io_dataOut_7_1_4(dataModule_io_dataOut_7_1_4),
    .io_dataOut_7_1_5(dataModule_io_dataOut_7_1_5),
    .io_dataOut_7_1_6(dataModule_io_dataOut_7_1_6),
    .io_dataOut_7_1_7(dataModule_io_dataOut_7_1_7),
    .io_dataOut_7_2_0(dataModule_io_dataOut_7_2_0),
    .io_dataOut_7_2_1(dataModule_io_dataOut_7_2_1),
    .io_dataOut_7_2_2(dataModule_io_dataOut_7_2_2),
    .io_dataOut_7_2_3(dataModule_io_dataOut_7_2_3),
    .io_dataOut_7_2_4(dataModule_io_dataOut_7_2_4),
    .io_dataOut_7_2_5(dataModule_io_dataOut_7_2_5),
    .io_dataOut_7_2_6(dataModule_io_dataOut_7_2_6),
    .io_dataOut_7_2_7(dataModule_io_dataOut_7_2_7),
    .io_dataOut_7_3_0(dataModule_io_dataOut_7_3_0),
    .io_dataOut_7_3_1(dataModule_io_dataOut_7_3_1),
    .io_dataOut_7_3_2(dataModule_io_dataOut_7_3_2),
    .io_dataOut_7_3_3(dataModule_io_dataOut_7_3_3),
    .io_dataOut_7_3_4(dataModule_io_dataOut_7_3_4),
    .io_dataOut_7_3_5(dataModule_io_dataOut_7_3_5),
    .io_dataOut_7_3_6(dataModule_io_dataOut_7_3_6),
    .io_dataOut_7_3_7(dataModule_io_dataOut_7_3_7),
    .io_dataOut_7_4_0(dataModule_io_dataOut_7_4_0),
    .io_dataOut_7_4_1(dataModule_io_dataOut_7_4_1),
    .io_dataOut_7_4_2(dataModule_io_dataOut_7_4_2),
    .io_dataOut_7_4_3(dataModule_io_dataOut_7_4_3),
    .io_dataOut_7_4_4(dataModule_io_dataOut_7_4_4),
    .io_dataOut_7_4_5(dataModule_io_dataOut_7_4_5),
    .io_dataOut_7_4_6(dataModule_io_dataOut_7_4_6),
    .io_dataOut_7_4_7(dataModule_io_dataOut_7_4_7),
    .io_dataOut_7_5_0(dataModule_io_dataOut_7_5_0),
    .io_dataOut_7_5_1(dataModule_io_dataOut_7_5_1),
    .io_dataOut_7_5_2(dataModule_io_dataOut_7_5_2),
    .io_dataOut_7_5_3(dataModule_io_dataOut_7_5_3),
    .io_dataOut_7_5_4(dataModule_io_dataOut_7_5_4),
    .io_dataOut_7_5_5(dataModule_io_dataOut_7_5_5),
    .io_dataOut_7_5_6(dataModule_io_dataOut_7_5_6),
    .io_dataOut_7_5_7(dataModule_io_dataOut_7_5_7),
    .io_dataOut_7_6_0(dataModule_io_dataOut_7_6_0),
    .io_dataOut_7_6_1(dataModule_io_dataOut_7_6_1),
    .io_dataOut_7_6_2(dataModule_io_dataOut_7_6_2),
    .io_dataOut_7_6_3(dataModule_io_dataOut_7_6_3),
    .io_dataOut_7_6_4(dataModule_io_dataOut_7_6_4),
    .io_dataOut_7_6_5(dataModule_io_dataOut_7_6_5),
    .io_dataOut_7_6_6(dataModule_io_dataOut_7_6_6),
    .io_dataOut_7_6_7(dataModule_io_dataOut_7_6_7),
    .io_dataOut_7_7_0(dataModule_io_dataOut_7_7_0),
    .io_dataOut_7_7_1(dataModule_io_dataOut_7_7_1),
    .io_dataOut_7_7_2(dataModule_io_dataOut_7_7_2),
    .io_dataOut_7_7_3(dataModule_io_dataOut_7_7_3),
    .io_dataOut_7_7_4(dataModule_io_dataOut_7_7_4),
    .io_dataOut_7_7_5(dataModule_io_dataOut_7_7_5),
    .io_dataOut_7_7_6(dataModule_io_dataOut_7_7_6),
    .io_dataOut_7_7_7(dataModule_io_dataOut_7_7_7),
    .io_dataOut_8_0_0(dataModule_io_dataOut_8_0_0),
    .io_dataOut_8_0_1(dataModule_io_dataOut_8_0_1),
    .io_dataOut_8_0_2(dataModule_io_dataOut_8_0_2),
    .io_dataOut_8_0_3(dataModule_io_dataOut_8_0_3),
    .io_dataOut_8_0_4(dataModule_io_dataOut_8_0_4),
    .io_dataOut_8_0_5(dataModule_io_dataOut_8_0_5),
    .io_dataOut_8_0_6(dataModule_io_dataOut_8_0_6),
    .io_dataOut_8_0_7(dataModule_io_dataOut_8_0_7),
    .io_dataOut_8_1_0(dataModule_io_dataOut_8_1_0),
    .io_dataOut_8_1_1(dataModule_io_dataOut_8_1_1),
    .io_dataOut_8_1_2(dataModule_io_dataOut_8_1_2),
    .io_dataOut_8_1_3(dataModule_io_dataOut_8_1_3),
    .io_dataOut_8_1_4(dataModule_io_dataOut_8_1_4),
    .io_dataOut_8_1_5(dataModule_io_dataOut_8_1_5),
    .io_dataOut_8_1_6(dataModule_io_dataOut_8_1_6),
    .io_dataOut_8_1_7(dataModule_io_dataOut_8_1_7),
    .io_dataOut_8_2_0(dataModule_io_dataOut_8_2_0),
    .io_dataOut_8_2_1(dataModule_io_dataOut_8_2_1),
    .io_dataOut_8_2_2(dataModule_io_dataOut_8_2_2),
    .io_dataOut_8_2_3(dataModule_io_dataOut_8_2_3),
    .io_dataOut_8_2_4(dataModule_io_dataOut_8_2_4),
    .io_dataOut_8_2_5(dataModule_io_dataOut_8_2_5),
    .io_dataOut_8_2_6(dataModule_io_dataOut_8_2_6),
    .io_dataOut_8_2_7(dataModule_io_dataOut_8_2_7),
    .io_dataOut_8_3_0(dataModule_io_dataOut_8_3_0),
    .io_dataOut_8_3_1(dataModule_io_dataOut_8_3_1),
    .io_dataOut_8_3_2(dataModule_io_dataOut_8_3_2),
    .io_dataOut_8_3_3(dataModule_io_dataOut_8_3_3),
    .io_dataOut_8_3_4(dataModule_io_dataOut_8_3_4),
    .io_dataOut_8_3_5(dataModule_io_dataOut_8_3_5),
    .io_dataOut_8_3_6(dataModule_io_dataOut_8_3_6),
    .io_dataOut_8_3_7(dataModule_io_dataOut_8_3_7),
    .io_dataOut_8_4_0(dataModule_io_dataOut_8_4_0),
    .io_dataOut_8_4_1(dataModule_io_dataOut_8_4_1),
    .io_dataOut_8_4_2(dataModule_io_dataOut_8_4_2),
    .io_dataOut_8_4_3(dataModule_io_dataOut_8_4_3),
    .io_dataOut_8_4_4(dataModule_io_dataOut_8_4_4),
    .io_dataOut_8_4_5(dataModule_io_dataOut_8_4_5),
    .io_dataOut_8_4_6(dataModule_io_dataOut_8_4_6),
    .io_dataOut_8_4_7(dataModule_io_dataOut_8_4_7),
    .io_dataOut_8_5_0(dataModule_io_dataOut_8_5_0),
    .io_dataOut_8_5_1(dataModule_io_dataOut_8_5_1),
    .io_dataOut_8_5_2(dataModule_io_dataOut_8_5_2),
    .io_dataOut_8_5_3(dataModule_io_dataOut_8_5_3),
    .io_dataOut_8_5_4(dataModule_io_dataOut_8_5_4),
    .io_dataOut_8_5_5(dataModule_io_dataOut_8_5_5),
    .io_dataOut_8_5_6(dataModule_io_dataOut_8_5_6),
    .io_dataOut_8_5_7(dataModule_io_dataOut_8_5_7),
    .io_dataOut_8_6_0(dataModule_io_dataOut_8_6_0),
    .io_dataOut_8_6_1(dataModule_io_dataOut_8_6_1),
    .io_dataOut_8_6_2(dataModule_io_dataOut_8_6_2),
    .io_dataOut_8_6_3(dataModule_io_dataOut_8_6_3),
    .io_dataOut_8_6_4(dataModule_io_dataOut_8_6_4),
    .io_dataOut_8_6_5(dataModule_io_dataOut_8_6_5),
    .io_dataOut_8_6_6(dataModule_io_dataOut_8_6_6),
    .io_dataOut_8_6_7(dataModule_io_dataOut_8_6_7),
    .io_dataOut_8_7_0(dataModule_io_dataOut_8_7_0),
    .io_dataOut_8_7_1(dataModule_io_dataOut_8_7_1),
    .io_dataOut_8_7_2(dataModule_io_dataOut_8_7_2),
    .io_dataOut_8_7_3(dataModule_io_dataOut_8_7_3),
    .io_dataOut_8_7_4(dataModule_io_dataOut_8_7_4),
    .io_dataOut_8_7_5(dataModule_io_dataOut_8_7_5),
    .io_dataOut_8_7_6(dataModule_io_dataOut_8_7_6),
    .io_dataOut_8_7_7(dataModule_io_dataOut_8_7_7),
    .io_dataOut_9_0_0(dataModule_io_dataOut_9_0_0),
    .io_dataOut_9_0_1(dataModule_io_dataOut_9_0_1),
    .io_dataOut_9_0_2(dataModule_io_dataOut_9_0_2),
    .io_dataOut_9_0_3(dataModule_io_dataOut_9_0_3),
    .io_dataOut_9_0_4(dataModule_io_dataOut_9_0_4),
    .io_dataOut_9_0_5(dataModule_io_dataOut_9_0_5),
    .io_dataOut_9_0_6(dataModule_io_dataOut_9_0_6),
    .io_dataOut_9_0_7(dataModule_io_dataOut_9_0_7),
    .io_dataOut_9_1_0(dataModule_io_dataOut_9_1_0),
    .io_dataOut_9_1_1(dataModule_io_dataOut_9_1_1),
    .io_dataOut_9_1_2(dataModule_io_dataOut_9_1_2),
    .io_dataOut_9_1_3(dataModule_io_dataOut_9_1_3),
    .io_dataOut_9_1_4(dataModule_io_dataOut_9_1_4),
    .io_dataOut_9_1_5(dataModule_io_dataOut_9_1_5),
    .io_dataOut_9_1_6(dataModule_io_dataOut_9_1_6),
    .io_dataOut_9_1_7(dataModule_io_dataOut_9_1_7),
    .io_dataOut_9_2_0(dataModule_io_dataOut_9_2_0),
    .io_dataOut_9_2_1(dataModule_io_dataOut_9_2_1),
    .io_dataOut_9_2_2(dataModule_io_dataOut_9_2_2),
    .io_dataOut_9_2_3(dataModule_io_dataOut_9_2_3),
    .io_dataOut_9_2_4(dataModule_io_dataOut_9_2_4),
    .io_dataOut_9_2_5(dataModule_io_dataOut_9_2_5),
    .io_dataOut_9_2_6(dataModule_io_dataOut_9_2_6),
    .io_dataOut_9_2_7(dataModule_io_dataOut_9_2_7),
    .io_dataOut_9_3_0(dataModule_io_dataOut_9_3_0),
    .io_dataOut_9_3_1(dataModule_io_dataOut_9_3_1),
    .io_dataOut_9_3_2(dataModule_io_dataOut_9_3_2),
    .io_dataOut_9_3_3(dataModule_io_dataOut_9_3_3),
    .io_dataOut_9_3_4(dataModule_io_dataOut_9_3_4),
    .io_dataOut_9_3_5(dataModule_io_dataOut_9_3_5),
    .io_dataOut_9_3_6(dataModule_io_dataOut_9_3_6),
    .io_dataOut_9_3_7(dataModule_io_dataOut_9_3_7),
    .io_dataOut_9_4_0(dataModule_io_dataOut_9_4_0),
    .io_dataOut_9_4_1(dataModule_io_dataOut_9_4_1),
    .io_dataOut_9_4_2(dataModule_io_dataOut_9_4_2),
    .io_dataOut_9_4_3(dataModule_io_dataOut_9_4_3),
    .io_dataOut_9_4_4(dataModule_io_dataOut_9_4_4),
    .io_dataOut_9_4_5(dataModule_io_dataOut_9_4_5),
    .io_dataOut_9_4_6(dataModule_io_dataOut_9_4_6),
    .io_dataOut_9_4_7(dataModule_io_dataOut_9_4_7),
    .io_dataOut_9_5_0(dataModule_io_dataOut_9_5_0),
    .io_dataOut_9_5_1(dataModule_io_dataOut_9_5_1),
    .io_dataOut_9_5_2(dataModule_io_dataOut_9_5_2),
    .io_dataOut_9_5_3(dataModule_io_dataOut_9_5_3),
    .io_dataOut_9_5_4(dataModule_io_dataOut_9_5_4),
    .io_dataOut_9_5_5(dataModule_io_dataOut_9_5_5),
    .io_dataOut_9_5_6(dataModule_io_dataOut_9_5_6),
    .io_dataOut_9_5_7(dataModule_io_dataOut_9_5_7),
    .io_dataOut_9_6_0(dataModule_io_dataOut_9_6_0),
    .io_dataOut_9_6_1(dataModule_io_dataOut_9_6_1),
    .io_dataOut_9_6_2(dataModule_io_dataOut_9_6_2),
    .io_dataOut_9_6_3(dataModule_io_dataOut_9_6_3),
    .io_dataOut_9_6_4(dataModule_io_dataOut_9_6_4),
    .io_dataOut_9_6_5(dataModule_io_dataOut_9_6_5),
    .io_dataOut_9_6_6(dataModule_io_dataOut_9_6_6),
    .io_dataOut_9_6_7(dataModule_io_dataOut_9_6_7),
    .io_dataOut_9_7_0(dataModule_io_dataOut_9_7_0),
    .io_dataOut_9_7_1(dataModule_io_dataOut_9_7_1),
    .io_dataOut_9_7_2(dataModule_io_dataOut_9_7_2),
    .io_dataOut_9_7_3(dataModule_io_dataOut_9_7_3),
    .io_dataOut_9_7_4(dataModule_io_dataOut_9_7_4),
    .io_dataOut_9_7_5(dataModule_io_dataOut_9_7_5),
    .io_dataOut_9_7_6(dataModule_io_dataOut_9_7_6),
    .io_dataOut_9_7_7(dataModule_io_dataOut_9_7_7),
    .io_dataOut_10_0_0(dataModule_io_dataOut_10_0_0),
    .io_dataOut_10_0_1(dataModule_io_dataOut_10_0_1),
    .io_dataOut_10_0_2(dataModule_io_dataOut_10_0_2),
    .io_dataOut_10_0_3(dataModule_io_dataOut_10_0_3),
    .io_dataOut_10_0_4(dataModule_io_dataOut_10_0_4),
    .io_dataOut_10_0_5(dataModule_io_dataOut_10_0_5),
    .io_dataOut_10_0_6(dataModule_io_dataOut_10_0_6),
    .io_dataOut_10_0_7(dataModule_io_dataOut_10_0_7),
    .io_dataOut_10_1_0(dataModule_io_dataOut_10_1_0),
    .io_dataOut_10_1_1(dataModule_io_dataOut_10_1_1),
    .io_dataOut_10_1_2(dataModule_io_dataOut_10_1_2),
    .io_dataOut_10_1_3(dataModule_io_dataOut_10_1_3),
    .io_dataOut_10_1_4(dataModule_io_dataOut_10_1_4),
    .io_dataOut_10_1_5(dataModule_io_dataOut_10_1_5),
    .io_dataOut_10_1_6(dataModule_io_dataOut_10_1_6),
    .io_dataOut_10_1_7(dataModule_io_dataOut_10_1_7),
    .io_dataOut_10_2_0(dataModule_io_dataOut_10_2_0),
    .io_dataOut_10_2_1(dataModule_io_dataOut_10_2_1),
    .io_dataOut_10_2_2(dataModule_io_dataOut_10_2_2),
    .io_dataOut_10_2_3(dataModule_io_dataOut_10_2_3),
    .io_dataOut_10_2_4(dataModule_io_dataOut_10_2_4),
    .io_dataOut_10_2_5(dataModule_io_dataOut_10_2_5),
    .io_dataOut_10_2_6(dataModule_io_dataOut_10_2_6),
    .io_dataOut_10_2_7(dataModule_io_dataOut_10_2_7),
    .io_dataOut_10_3_0(dataModule_io_dataOut_10_3_0),
    .io_dataOut_10_3_1(dataModule_io_dataOut_10_3_1),
    .io_dataOut_10_3_2(dataModule_io_dataOut_10_3_2),
    .io_dataOut_10_3_3(dataModule_io_dataOut_10_3_3),
    .io_dataOut_10_3_4(dataModule_io_dataOut_10_3_4),
    .io_dataOut_10_3_5(dataModule_io_dataOut_10_3_5),
    .io_dataOut_10_3_6(dataModule_io_dataOut_10_3_6),
    .io_dataOut_10_3_7(dataModule_io_dataOut_10_3_7),
    .io_dataOut_10_4_0(dataModule_io_dataOut_10_4_0),
    .io_dataOut_10_4_1(dataModule_io_dataOut_10_4_1),
    .io_dataOut_10_4_2(dataModule_io_dataOut_10_4_2),
    .io_dataOut_10_4_3(dataModule_io_dataOut_10_4_3),
    .io_dataOut_10_4_4(dataModule_io_dataOut_10_4_4),
    .io_dataOut_10_4_5(dataModule_io_dataOut_10_4_5),
    .io_dataOut_10_4_6(dataModule_io_dataOut_10_4_6),
    .io_dataOut_10_4_7(dataModule_io_dataOut_10_4_7),
    .io_dataOut_10_5_0(dataModule_io_dataOut_10_5_0),
    .io_dataOut_10_5_1(dataModule_io_dataOut_10_5_1),
    .io_dataOut_10_5_2(dataModule_io_dataOut_10_5_2),
    .io_dataOut_10_5_3(dataModule_io_dataOut_10_5_3),
    .io_dataOut_10_5_4(dataModule_io_dataOut_10_5_4),
    .io_dataOut_10_5_5(dataModule_io_dataOut_10_5_5),
    .io_dataOut_10_5_6(dataModule_io_dataOut_10_5_6),
    .io_dataOut_10_5_7(dataModule_io_dataOut_10_5_7),
    .io_dataOut_10_6_0(dataModule_io_dataOut_10_6_0),
    .io_dataOut_10_6_1(dataModule_io_dataOut_10_6_1),
    .io_dataOut_10_6_2(dataModule_io_dataOut_10_6_2),
    .io_dataOut_10_6_3(dataModule_io_dataOut_10_6_3),
    .io_dataOut_10_6_4(dataModule_io_dataOut_10_6_4),
    .io_dataOut_10_6_5(dataModule_io_dataOut_10_6_5),
    .io_dataOut_10_6_6(dataModule_io_dataOut_10_6_6),
    .io_dataOut_10_6_7(dataModule_io_dataOut_10_6_7),
    .io_dataOut_10_7_0(dataModule_io_dataOut_10_7_0),
    .io_dataOut_10_7_1(dataModule_io_dataOut_10_7_1),
    .io_dataOut_10_7_2(dataModule_io_dataOut_10_7_2),
    .io_dataOut_10_7_3(dataModule_io_dataOut_10_7_3),
    .io_dataOut_10_7_4(dataModule_io_dataOut_10_7_4),
    .io_dataOut_10_7_5(dataModule_io_dataOut_10_7_5),
    .io_dataOut_10_7_6(dataModule_io_dataOut_10_7_6),
    .io_dataOut_10_7_7(dataModule_io_dataOut_10_7_7),
    .io_dataOut_11_0_0(dataModule_io_dataOut_11_0_0),
    .io_dataOut_11_0_1(dataModule_io_dataOut_11_0_1),
    .io_dataOut_11_0_2(dataModule_io_dataOut_11_0_2),
    .io_dataOut_11_0_3(dataModule_io_dataOut_11_0_3),
    .io_dataOut_11_0_4(dataModule_io_dataOut_11_0_4),
    .io_dataOut_11_0_5(dataModule_io_dataOut_11_0_5),
    .io_dataOut_11_0_6(dataModule_io_dataOut_11_0_6),
    .io_dataOut_11_0_7(dataModule_io_dataOut_11_0_7),
    .io_dataOut_11_1_0(dataModule_io_dataOut_11_1_0),
    .io_dataOut_11_1_1(dataModule_io_dataOut_11_1_1),
    .io_dataOut_11_1_2(dataModule_io_dataOut_11_1_2),
    .io_dataOut_11_1_3(dataModule_io_dataOut_11_1_3),
    .io_dataOut_11_1_4(dataModule_io_dataOut_11_1_4),
    .io_dataOut_11_1_5(dataModule_io_dataOut_11_1_5),
    .io_dataOut_11_1_6(dataModule_io_dataOut_11_1_6),
    .io_dataOut_11_1_7(dataModule_io_dataOut_11_1_7),
    .io_dataOut_11_2_0(dataModule_io_dataOut_11_2_0),
    .io_dataOut_11_2_1(dataModule_io_dataOut_11_2_1),
    .io_dataOut_11_2_2(dataModule_io_dataOut_11_2_2),
    .io_dataOut_11_2_3(dataModule_io_dataOut_11_2_3),
    .io_dataOut_11_2_4(dataModule_io_dataOut_11_2_4),
    .io_dataOut_11_2_5(dataModule_io_dataOut_11_2_5),
    .io_dataOut_11_2_6(dataModule_io_dataOut_11_2_6),
    .io_dataOut_11_2_7(dataModule_io_dataOut_11_2_7),
    .io_dataOut_11_3_0(dataModule_io_dataOut_11_3_0),
    .io_dataOut_11_3_1(dataModule_io_dataOut_11_3_1),
    .io_dataOut_11_3_2(dataModule_io_dataOut_11_3_2),
    .io_dataOut_11_3_3(dataModule_io_dataOut_11_3_3),
    .io_dataOut_11_3_4(dataModule_io_dataOut_11_3_4),
    .io_dataOut_11_3_5(dataModule_io_dataOut_11_3_5),
    .io_dataOut_11_3_6(dataModule_io_dataOut_11_3_6),
    .io_dataOut_11_3_7(dataModule_io_dataOut_11_3_7),
    .io_dataOut_11_4_0(dataModule_io_dataOut_11_4_0),
    .io_dataOut_11_4_1(dataModule_io_dataOut_11_4_1),
    .io_dataOut_11_4_2(dataModule_io_dataOut_11_4_2),
    .io_dataOut_11_4_3(dataModule_io_dataOut_11_4_3),
    .io_dataOut_11_4_4(dataModule_io_dataOut_11_4_4),
    .io_dataOut_11_4_5(dataModule_io_dataOut_11_4_5),
    .io_dataOut_11_4_6(dataModule_io_dataOut_11_4_6),
    .io_dataOut_11_4_7(dataModule_io_dataOut_11_4_7),
    .io_dataOut_11_5_0(dataModule_io_dataOut_11_5_0),
    .io_dataOut_11_5_1(dataModule_io_dataOut_11_5_1),
    .io_dataOut_11_5_2(dataModule_io_dataOut_11_5_2),
    .io_dataOut_11_5_3(dataModule_io_dataOut_11_5_3),
    .io_dataOut_11_5_4(dataModule_io_dataOut_11_5_4),
    .io_dataOut_11_5_5(dataModule_io_dataOut_11_5_5),
    .io_dataOut_11_5_6(dataModule_io_dataOut_11_5_6),
    .io_dataOut_11_5_7(dataModule_io_dataOut_11_5_7),
    .io_dataOut_11_6_0(dataModule_io_dataOut_11_6_0),
    .io_dataOut_11_6_1(dataModule_io_dataOut_11_6_1),
    .io_dataOut_11_6_2(dataModule_io_dataOut_11_6_2),
    .io_dataOut_11_6_3(dataModule_io_dataOut_11_6_3),
    .io_dataOut_11_6_4(dataModule_io_dataOut_11_6_4),
    .io_dataOut_11_6_5(dataModule_io_dataOut_11_6_5),
    .io_dataOut_11_6_6(dataModule_io_dataOut_11_6_6),
    .io_dataOut_11_6_7(dataModule_io_dataOut_11_6_7),
    .io_dataOut_11_7_0(dataModule_io_dataOut_11_7_0),
    .io_dataOut_11_7_1(dataModule_io_dataOut_11_7_1),
    .io_dataOut_11_7_2(dataModule_io_dataOut_11_7_2),
    .io_dataOut_11_7_3(dataModule_io_dataOut_11_7_3),
    .io_dataOut_11_7_4(dataModule_io_dataOut_11_7_4),
    .io_dataOut_11_7_5(dataModule_io_dataOut_11_7_5),
    .io_dataOut_11_7_6(dataModule_io_dataOut_11_7_6),
    .io_dataOut_11_7_7(dataModule_io_dataOut_11_7_7),
    .io_dataOut_12_0_0(dataModule_io_dataOut_12_0_0),
    .io_dataOut_12_0_1(dataModule_io_dataOut_12_0_1),
    .io_dataOut_12_0_2(dataModule_io_dataOut_12_0_2),
    .io_dataOut_12_0_3(dataModule_io_dataOut_12_0_3),
    .io_dataOut_12_0_4(dataModule_io_dataOut_12_0_4),
    .io_dataOut_12_0_5(dataModule_io_dataOut_12_0_5),
    .io_dataOut_12_0_6(dataModule_io_dataOut_12_0_6),
    .io_dataOut_12_0_7(dataModule_io_dataOut_12_0_7),
    .io_dataOut_12_1_0(dataModule_io_dataOut_12_1_0),
    .io_dataOut_12_1_1(dataModule_io_dataOut_12_1_1),
    .io_dataOut_12_1_2(dataModule_io_dataOut_12_1_2),
    .io_dataOut_12_1_3(dataModule_io_dataOut_12_1_3),
    .io_dataOut_12_1_4(dataModule_io_dataOut_12_1_4),
    .io_dataOut_12_1_5(dataModule_io_dataOut_12_1_5),
    .io_dataOut_12_1_6(dataModule_io_dataOut_12_1_6),
    .io_dataOut_12_1_7(dataModule_io_dataOut_12_1_7),
    .io_dataOut_12_2_0(dataModule_io_dataOut_12_2_0),
    .io_dataOut_12_2_1(dataModule_io_dataOut_12_2_1),
    .io_dataOut_12_2_2(dataModule_io_dataOut_12_2_2),
    .io_dataOut_12_2_3(dataModule_io_dataOut_12_2_3),
    .io_dataOut_12_2_4(dataModule_io_dataOut_12_2_4),
    .io_dataOut_12_2_5(dataModule_io_dataOut_12_2_5),
    .io_dataOut_12_2_6(dataModule_io_dataOut_12_2_6),
    .io_dataOut_12_2_7(dataModule_io_dataOut_12_2_7),
    .io_dataOut_12_3_0(dataModule_io_dataOut_12_3_0),
    .io_dataOut_12_3_1(dataModule_io_dataOut_12_3_1),
    .io_dataOut_12_3_2(dataModule_io_dataOut_12_3_2),
    .io_dataOut_12_3_3(dataModule_io_dataOut_12_3_3),
    .io_dataOut_12_3_4(dataModule_io_dataOut_12_3_4),
    .io_dataOut_12_3_5(dataModule_io_dataOut_12_3_5),
    .io_dataOut_12_3_6(dataModule_io_dataOut_12_3_6),
    .io_dataOut_12_3_7(dataModule_io_dataOut_12_3_7),
    .io_dataOut_12_4_0(dataModule_io_dataOut_12_4_0),
    .io_dataOut_12_4_1(dataModule_io_dataOut_12_4_1),
    .io_dataOut_12_4_2(dataModule_io_dataOut_12_4_2),
    .io_dataOut_12_4_3(dataModule_io_dataOut_12_4_3),
    .io_dataOut_12_4_4(dataModule_io_dataOut_12_4_4),
    .io_dataOut_12_4_5(dataModule_io_dataOut_12_4_5),
    .io_dataOut_12_4_6(dataModule_io_dataOut_12_4_6),
    .io_dataOut_12_4_7(dataModule_io_dataOut_12_4_7),
    .io_dataOut_12_5_0(dataModule_io_dataOut_12_5_0),
    .io_dataOut_12_5_1(dataModule_io_dataOut_12_5_1),
    .io_dataOut_12_5_2(dataModule_io_dataOut_12_5_2),
    .io_dataOut_12_5_3(dataModule_io_dataOut_12_5_3),
    .io_dataOut_12_5_4(dataModule_io_dataOut_12_5_4),
    .io_dataOut_12_5_5(dataModule_io_dataOut_12_5_5),
    .io_dataOut_12_5_6(dataModule_io_dataOut_12_5_6),
    .io_dataOut_12_5_7(dataModule_io_dataOut_12_5_7),
    .io_dataOut_12_6_0(dataModule_io_dataOut_12_6_0),
    .io_dataOut_12_6_1(dataModule_io_dataOut_12_6_1),
    .io_dataOut_12_6_2(dataModule_io_dataOut_12_6_2),
    .io_dataOut_12_6_3(dataModule_io_dataOut_12_6_3),
    .io_dataOut_12_6_4(dataModule_io_dataOut_12_6_4),
    .io_dataOut_12_6_5(dataModule_io_dataOut_12_6_5),
    .io_dataOut_12_6_6(dataModule_io_dataOut_12_6_6),
    .io_dataOut_12_6_7(dataModule_io_dataOut_12_6_7),
    .io_dataOut_12_7_0(dataModule_io_dataOut_12_7_0),
    .io_dataOut_12_7_1(dataModule_io_dataOut_12_7_1),
    .io_dataOut_12_7_2(dataModule_io_dataOut_12_7_2),
    .io_dataOut_12_7_3(dataModule_io_dataOut_12_7_3),
    .io_dataOut_12_7_4(dataModule_io_dataOut_12_7_4),
    .io_dataOut_12_7_5(dataModule_io_dataOut_12_7_5),
    .io_dataOut_12_7_6(dataModule_io_dataOut_12_7_6),
    .io_dataOut_12_7_7(dataModule_io_dataOut_12_7_7),
    .io_dataOut_13_0_0(dataModule_io_dataOut_13_0_0),
    .io_dataOut_13_0_1(dataModule_io_dataOut_13_0_1),
    .io_dataOut_13_0_2(dataModule_io_dataOut_13_0_2),
    .io_dataOut_13_0_3(dataModule_io_dataOut_13_0_3),
    .io_dataOut_13_0_4(dataModule_io_dataOut_13_0_4),
    .io_dataOut_13_0_5(dataModule_io_dataOut_13_0_5),
    .io_dataOut_13_0_6(dataModule_io_dataOut_13_0_6),
    .io_dataOut_13_0_7(dataModule_io_dataOut_13_0_7),
    .io_dataOut_13_1_0(dataModule_io_dataOut_13_1_0),
    .io_dataOut_13_1_1(dataModule_io_dataOut_13_1_1),
    .io_dataOut_13_1_2(dataModule_io_dataOut_13_1_2),
    .io_dataOut_13_1_3(dataModule_io_dataOut_13_1_3),
    .io_dataOut_13_1_4(dataModule_io_dataOut_13_1_4),
    .io_dataOut_13_1_5(dataModule_io_dataOut_13_1_5),
    .io_dataOut_13_1_6(dataModule_io_dataOut_13_1_6),
    .io_dataOut_13_1_7(dataModule_io_dataOut_13_1_7),
    .io_dataOut_13_2_0(dataModule_io_dataOut_13_2_0),
    .io_dataOut_13_2_1(dataModule_io_dataOut_13_2_1),
    .io_dataOut_13_2_2(dataModule_io_dataOut_13_2_2),
    .io_dataOut_13_2_3(dataModule_io_dataOut_13_2_3),
    .io_dataOut_13_2_4(dataModule_io_dataOut_13_2_4),
    .io_dataOut_13_2_5(dataModule_io_dataOut_13_2_5),
    .io_dataOut_13_2_6(dataModule_io_dataOut_13_2_6),
    .io_dataOut_13_2_7(dataModule_io_dataOut_13_2_7),
    .io_dataOut_13_3_0(dataModule_io_dataOut_13_3_0),
    .io_dataOut_13_3_1(dataModule_io_dataOut_13_3_1),
    .io_dataOut_13_3_2(dataModule_io_dataOut_13_3_2),
    .io_dataOut_13_3_3(dataModule_io_dataOut_13_3_3),
    .io_dataOut_13_3_4(dataModule_io_dataOut_13_3_4),
    .io_dataOut_13_3_5(dataModule_io_dataOut_13_3_5),
    .io_dataOut_13_3_6(dataModule_io_dataOut_13_3_6),
    .io_dataOut_13_3_7(dataModule_io_dataOut_13_3_7),
    .io_dataOut_13_4_0(dataModule_io_dataOut_13_4_0),
    .io_dataOut_13_4_1(dataModule_io_dataOut_13_4_1),
    .io_dataOut_13_4_2(dataModule_io_dataOut_13_4_2),
    .io_dataOut_13_4_3(dataModule_io_dataOut_13_4_3),
    .io_dataOut_13_4_4(dataModule_io_dataOut_13_4_4),
    .io_dataOut_13_4_5(dataModule_io_dataOut_13_4_5),
    .io_dataOut_13_4_6(dataModule_io_dataOut_13_4_6),
    .io_dataOut_13_4_7(dataModule_io_dataOut_13_4_7),
    .io_dataOut_13_5_0(dataModule_io_dataOut_13_5_0),
    .io_dataOut_13_5_1(dataModule_io_dataOut_13_5_1),
    .io_dataOut_13_5_2(dataModule_io_dataOut_13_5_2),
    .io_dataOut_13_5_3(dataModule_io_dataOut_13_5_3),
    .io_dataOut_13_5_4(dataModule_io_dataOut_13_5_4),
    .io_dataOut_13_5_5(dataModule_io_dataOut_13_5_5),
    .io_dataOut_13_5_6(dataModule_io_dataOut_13_5_6),
    .io_dataOut_13_5_7(dataModule_io_dataOut_13_5_7),
    .io_dataOut_13_6_0(dataModule_io_dataOut_13_6_0),
    .io_dataOut_13_6_1(dataModule_io_dataOut_13_6_1),
    .io_dataOut_13_6_2(dataModule_io_dataOut_13_6_2),
    .io_dataOut_13_6_3(dataModule_io_dataOut_13_6_3),
    .io_dataOut_13_6_4(dataModule_io_dataOut_13_6_4),
    .io_dataOut_13_6_5(dataModule_io_dataOut_13_6_5),
    .io_dataOut_13_6_6(dataModule_io_dataOut_13_6_6),
    .io_dataOut_13_6_7(dataModule_io_dataOut_13_6_7),
    .io_dataOut_13_7_0(dataModule_io_dataOut_13_7_0),
    .io_dataOut_13_7_1(dataModule_io_dataOut_13_7_1),
    .io_dataOut_13_7_2(dataModule_io_dataOut_13_7_2),
    .io_dataOut_13_7_3(dataModule_io_dataOut_13_7_3),
    .io_dataOut_13_7_4(dataModule_io_dataOut_13_7_4),
    .io_dataOut_13_7_5(dataModule_io_dataOut_13_7_5),
    .io_dataOut_13_7_6(dataModule_io_dataOut_13_7_6),
    .io_dataOut_13_7_7(dataModule_io_dataOut_13_7_7),
    .io_dataOut_14_0_0(dataModule_io_dataOut_14_0_0),
    .io_dataOut_14_0_1(dataModule_io_dataOut_14_0_1),
    .io_dataOut_14_0_2(dataModule_io_dataOut_14_0_2),
    .io_dataOut_14_0_3(dataModule_io_dataOut_14_0_3),
    .io_dataOut_14_0_4(dataModule_io_dataOut_14_0_4),
    .io_dataOut_14_0_5(dataModule_io_dataOut_14_0_5),
    .io_dataOut_14_0_6(dataModule_io_dataOut_14_0_6),
    .io_dataOut_14_0_7(dataModule_io_dataOut_14_0_7),
    .io_dataOut_14_1_0(dataModule_io_dataOut_14_1_0),
    .io_dataOut_14_1_1(dataModule_io_dataOut_14_1_1),
    .io_dataOut_14_1_2(dataModule_io_dataOut_14_1_2),
    .io_dataOut_14_1_3(dataModule_io_dataOut_14_1_3),
    .io_dataOut_14_1_4(dataModule_io_dataOut_14_1_4),
    .io_dataOut_14_1_5(dataModule_io_dataOut_14_1_5),
    .io_dataOut_14_1_6(dataModule_io_dataOut_14_1_6),
    .io_dataOut_14_1_7(dataModule_io_dataOut_14_1_7),
    .io_dataOut_14_2_0(dataModule_io_dataOut_14_2_0),
    .io_dataOut_14_2_1(dataModule_io_dataOut_14_2_1),
    .io_dataOut_14_2_2(dataModule_io_dataOut_14_2_2),
    .io_dataOut_14_2_3(dataModule_io_dataOut_14_2_3),
    .io_dataOut_14_2_4(dataModule_io_dataOut_14_2_4),
    .io_dataOut_14_2_5(dataModule_io_dataOut_14_2_5),
    .io_dataOut_14_2_6(dataModule_io_dataOut_14_2_6),
    .io_dataOut_14_2_7(dataModule_io_dataOut_14_2_7),
    .io_dataOut_14_3_0(dataModule_io_dataOut_14_3_0),
    .io_dataOut_14_3_1(dataModule_io_dataOut_14_3_1),
    .io_dataOut_14_3_2(dataModule_io_dataOut_14_3_2),
    .io_dataOut_14_3_3(dataModule_io_dataOut_14_3_3),
    .io_dataOut_14_3_4(dataModule_io_dataOut_14_3_4),
    .io_dataOut_14_3_5(dataModule_io_dataOut_14_3_5),
    .io_dataOut_14_3_6(dataModule_io_dataOut_14_3_6),
    .io_dataOut_14_3_7(dataModule_io_dataOut_14_3_7),
    .io_dataOut_14_4_0(dataModule_io_dataOut_14_4_0),
    .io_dataOut_14_4_1(dataModule_io_dataOut_14_4_1),
    .io_dataOut_14_4_2(dataModule_io_dataOut_14_4_2),
    .io_dataOut_14_4_3(dataModule_io_dataOut_14_4_3),
    .io_dataOut_14_4_4(dataModule_io_dataOut_14_4_4),
    .io_dataOut_14_4_5(dataModule_io_dataOut_14_4_5),
    .io_dataOut_14_4_6(dataModule_io_dataOut_14_4_6),
    .io_dataOut_14_4_7(dataModule_io_dataOut_14_4_7),
    .io_dataOut_14_5_0(dataModule_io_dataOut_14_5_0),
    .io_dataOut_14_5_1(dataModule_io_dataOut_14_5_1),
    .io_dataOut_14_5_2(dataModule_io_dataOut_14_5_2),
    .io_dataOut_14_5_3(dataModule_io_dataOut_14_5_3),
    .io_dataOut_14_5_4(dataModule_io_dataOut_14_5_4),
    .io_dataOut_14_5_5(dataModule_io_dataOut_14_5_5),
    .io_dataOut_14_5_6(dataModule_io_dataOut_14_5_6),
    .io_dataOut_14_5_7(dataModule_io_dataOut_14_5_7),
    .io_dataOut_14_6_0(dataModule_io_dataOut_14_6_0),
    .io_dataOut_14_6_1(dataModule_io_dataOut_14_6_1),
    .io_dataOut_14_6_2(dataModule_io_dataOut_14_6_2),
    .io_dataOut_14_6_3(dataModule_io_dataOut_14_6_3),
    .io_dataOut_14_6_4(dataModule_io_dataOut_14_6_4),
    .io_dataOut_14_6_5(dataModule_io_dataOut_14_6_5),
    .io_dataOut_14_6_6(dataModule_io_dataOut_14_6_6),
    .io_dataOut_14_6_7(dataModule_io_dataOut_14_6_7),
    .io_dataOut_14_7_0(dataModule_io_dataOut_14_7_0),
    .io_dataOut_14_7_1(dataModule_io_dataOut_14_7_1),
    .io_dataOut_14_7_2(dataModule_io_dataOut_14_7_2),
    .io_dataOut_14_7_3(dataModule_io_dataOut_14_7_3),
    .io_dataOut_14_7_4(dataModule_io_dataOut_14_7_4),
    .io_dataOut_14_7_5(dataModule_io_dataOut_14_7_5),
    .io_dataOut_14_7_6(dataModule_io_dataOut_14_7_6),
    .io_dataOut_14_7_7(dataModule_io_dataOut_14_7_7),
    .io_dataOut_15_0_0(dataModule_io_dataOut_15_0_0),
    .io_dataOut_15_0_1(dataModule_io_dataOut_15_0_1),
    .io_dataOut_15_0_2(dataModule_io_dataOut_15_0_2),
    .io_dataOut_15_0_3(dataModule_io_dataOut_15_0_3),
    .io_dataOut_15_0_4(dataModule_io_dataOut_15_0_4),
    .io_dataOut_15_0_5(dataModule_io_dataOut_15_0_5),
    .io_dataOut_15_0_6(dataModule_io_dataOut_15_0_6),
    .io_dataOut_15_0_7(dataModule_io_dataOut_15_0_7),
    .io_dataOut_15_1_0(dataModule_io_dataOut_15_1_0),
    .io_dataOut_15_1_1(dataModule_io_dataOut_15_1_1),
    .io_dataOut_15_1_2(dataModule_io_dataOut_15_1_2),
    .io_dataOut_15_1_3(dataModule_io_dataOut_15_1_3),
    .io_dataOut_15_1_4(dataModule_io_dataOut_15_1_4),
    .io_dataOut_15_1_5(dataModule_io_dataOut_15_1_5),
    .io_dataOut_15_1_6(dataModule_io_dataOut_15_1_6),
    .io_dataOut_15_1_7(dataModule_io_dataOut_15_1_7),
    .io_dataOut_15_2_0(dataModule_io_dataOut_15_2_0),
    .io_dataOut_15_2_1(dataModule_io_dataOut_15_2_1),
    .io_dataOut_15_2_2(dataModule_io_dataOut_15_2_2),
    .io_dataOut_15_2_3(dataModule_io_dataOut_15_2_3),
    .io_dataOut_15_2_4(dataModule_io_dataOut_15_2_4),
    .io_dataOut_15_2_5(dataModule_io_dataOut_15_2_5),
    .io_dataOut_15_2_6(dataModule_io_dataOut_15_2_6),
    .io_dataOut_15_2_7(dataModule_io_dataOut_15_2_7),
    .io_dataOut_15_3_0(dataModule_io_dataOut_15_3_0),
    .io_dataOut_15_3_1(dataModule_io_dataOut_15_3_1),
    .io_dataOut_15_3_2(dataModule_io_dataOut_15_3_2),
    .io_dataOut_15_3_3(dataModule_io_dataOut_15_3_3),
    .io_dataOut_15_3_4(dataModule_io_dataOut_15_3_4),
    .io_dataOut_15_3_5(dataModule_io_dataOut_15_3_5),
    .io_dataOut_15_3_6(dataModule_io_dataOut_15_3_6),
    .io_dataOut_15_3_7(dataModule_io_dataOut_15_3_7),
    .io_dataOut_15_4_0(dataModule_io_dataOut_15_4_0),
    .io_dataOut_15_4_1(dataModule_io_dataOut_15_4_1),
    .io_dataOut_15_4_2(dataModule_io_dataOut_15_4_2),
    .io_dataOut_15_4_3(dataModule_io_dataOut_15_4_3),
    .io_dataOut_15_4_4(dataModule_io_dataOut_15_4_4),
    .io_dataOut_15_4_5(dataModule_io_dataOut_15_4_5),
    .io_dataOut_15_4_6(dataModule_io_dataOut_15_4_6),
    .io_dataOut_15_4_7(dataModule_io_dataOut_15_4_7),
    .io_dataOut_15_5_0(dataModule_io_dataOut_15_5_0),
    .io_dataOut_15_5_1(dataModule_io_dataOut_15_5_1),
    .io_dataOut_15_5_2(dataModule_io_dataOut_15_5_2),
    .io_dataOut_15_5_3(dataModule_io_dataOut_15_5_3),
    .io_dataOut_15_5_4(dataModule_io_dataOut_15_5_4),
    .io_dataOut_15_5_5(dataModule_io_dataOut_15_5_5),
    .io_dataOut_15_5_6(dataModule_io_dataOut_15_5_6),
    .io_dataOut_15_5_7(dataModule_io_dataOut_15_5_7),
    .io_dataOut_15_6_0(dataModule_io_dataOut_15_6_0),
    .io_dataOut_15_6_1(dataModule_io_dataOut_15_6_1),
    .io_dataOut_15_6_2(dataModule_io_dataOut_15_6_2),
    .io_dataOut_15_6_3(dataModule_io_dataOut_15_6_3),
    .io_dataOut_15_6_4(dataModule_io_dataOut_15_6_4),
    .io_dataOut_15_6_5(dataModule_io_dataOut_15_6_5),
    .io_dataOut_15_6_6(dataModule_io_dataOut_15_6_6),
    .io_dataOut_15_6_7(dataModule_io_dataOut_15_6_7),
    .io_dataOut_15_7_0(dataModule_io_dataOut_15_7_0),
    .io_dataOut_15_7_1(dataModule_io_dataOut_15_7_1),
    .io_dataOut_15_7_2(dataModule_io_dataOut_15_7_2),
    .io_dataOut_15_7_3(dataModule_io_dataOut_15_7_3),
    .io_dataOut_15_7_4(dataModule_io_dataOut_15_7_4),
    .io_dataOut_15_7_5(dataModule_io_dataOut_15_7_5),
    .io_dataOut_15_7_6(dataModule_io_dataOut_15_7_6),
    .io_dataOut_15_7_7(dataModule_io_dataOut_15_7_7),
    .io_maskOut_0_0_0(dataModule_io_maskOut_0_0_0),
    .io_maskOut_0_0_1(dataModule_io_maskOut_0_0_1),
    .io_maskOut_0_0_2(dataModule_io_maskOut_0_0_2),
    .io_maskOut_0_0_3(dataModule_io_maskOut_0_0_3),
    .io_maskOut_0_0_4(dataModule_io_maskOut_0_0_4),
    .io_maskOut_0_0_5(dataModule_io_maskOut_0_0_5),
    .io_maskOut_0_0_6(dataModule_io_maskOut_0_0_6),
    .io_maskOut_0_0_7(dataModule_io_maskOut_0_0_7),
    .io_maskOut_0_1_0(dataModule_io_maskOut_0_1_0),
    .io_maskOut_0_1_1(dataModule_io_maskOut_0_1_1),
    .io_maskOut_0_1_2(dataModule_io_maskOut_0_1_2),
    .io_maskOut_0_1_3(dataModule_io_maskOut_0_1_3),
    .io_maskOut_0_1_4(dataModule_io_maskOut_0_1_4),
    .io_maskOut_0_1_5(dataModule_io_maskOut_0_1_5),
    .io_maskOut_0_1_6(dataModule_io_maskOut_0_1_6),
    .io_maskOut_0_1_7(dataModule_io_maskOut_0_1_7),
    .io_maskOut_0_2_0(dataModule_io_maskOut_0_2_0),
    .io_maskOut_0_2_1(dataModule_io_maskOut_0_2_1),
    .io_maskOut_0_2_2(dataModule_io_maskOut_0_2_2),
    .io_maskOut_0_2_3(dataModule_io_maskOut_0_2_3),
    .io_maskOut_0_2_4(dataModule_io_maskOut_0_2_4),
    .io_maskOut_0_2_5(dataModule_io_maskOut_0_2_5),
    .io_maskOut_0_2_6(dataModule_io_maskOut_0_2_6),
    .io_maskOut_0_2_7(dataModule_io_maskOut_0_2_7),
    .io_maskOut_0_3_0(dataModule_io_maskOut_0_3_0),
    .io_maskOut_0_3_1(dataModule_io_maskOut_0_3_1),
    .io_maskOut_0_3_2(dataModule_io_maskOut_0_3_2),
    .io_maskOut_0_3_3(dataModule_io_maskOut_0_3_3),
    .io_maskOut_0_3_4(dataModule_io_maskOut_0_3_4),
    .io_maskOut_0_3_5(dataModule_io_maskOut_0_3_5),
    .io_maskOut_0_3_6(dataModule_io_maskOut_0_3_6),
    .io_maskOut_0_3_7(dataModule_io_maskOut_0_3_7),
    .io_maskOut_0_4_0(dataModule_io_maskOut_0_4_0),
    .io_maskOut_0_4_1(dataModule_io_maskOut_0_4_1),
    .io_maskOut_0_4_2(dataModule_io_maskOut_0_4_2),
    .io_maskOut_0_4_3(dataModule_io_maskOut_0_4_3),
    .io_maskOut_0_4_4(dataModule_io_maskOut_0_4_4),
    .io_maskOut_0_4_5(dataModule_io_maskOut_0_4_5),
    .io_maskOut_0_4_6(dataModule_io_maskOut_0_4_6),
    .io_maskOut_0_4_7(dataModule_io_maskOut_0_4_7),
    .io_maskOut_0_5_0(dataModule_io_maskOut_0_5_0),
    .io_maskOut_0_5_1(dataModule_io_maskOut_0_5_1),
    .io_maskOut_0_5_2(dataModule_io_maskOut_0_5_2),
    .io_maskOut_0_5_3(dataModule_io_maskOut_0_5_3),
    .io_maskOut_0_5_4(dataModule_io_maskOut_0_5_4),
    .io_maskOut_0_5_5(dataModule_io_maskOut_0_5_5),
    .io_maskOut_0_5_6(dataModule_io_maskOut_0_5_6),
    .io_maskOut_0_5_7(dataModule_io_maskOut_0_5_7),
    .io_maskOut_0_6_0(dataModule_io_maskOut_0_6_0),
    .io_maskOut_0_6_1(dataModule_io_maskOut_0_6_1),
    .io_maskOut_0_6_2(dataModule_io_maskOut_0_6_2),
    .io_maskOut_0_6_3(dataModule_io_maskOut_0_6_3),
    .io_maskOut_0_6_4(dataModule_io_maskOut_0_6_4),
    .io_maskOut_0_6_5(dataModule_io_maskOut_0_6_5),
    .io_maskOut_0_6_6(dataModule_io_maskOut_0_6_6),
    .io_maskOut_0_6_7(dataModule_io_maskOut_0_6_7),
    .io_maskOut_0_7_0(dataModule_io_maskOut_0_7_0),
    .io_maskOut_0_7_1(dataModule_io_maskOut_0_7_1),
    .io_maskOut_0_7_2(dataModule_io_maskOut_0_7_2),
    .io_maskOut_0_7_3(dataModule_io_maskOut_0_7_3),
    .io_maskOut_0_7_4(dataModule_io_maskOut_0_7_4),
    .io_maskOut_0_7_5(dataModule_io_maskOut_0_7_5),
    .io_maskOut_0_7_6(dataModule_io_maskOut_0_7_6),
    .io_maskOut_0_7_7(dataModule_io_maskOut_0_7_7),
    .io_maskOut_1_0_0(dataModule_io_maskOut_1_0_0),
    .io_maskOut_1_0_1(dataModule_io_maskOut_1_0_1),
    .io_maskOut_1_0_2(dataModule_io_maskOut_1_0_2),
    .io_maskOut_1_0_3(dataModule_io_maskOut_1_0_3),
    .io_maskOut_1_0_4(dataModule_io_maskOut_1_0_4),
    .io_maskOut_1_0_5(dataModule_io_maskOut_1_0_5),
    .io_maskOut_1_0_6(dataModule_io_maskOut_1_0_6),
    .io_maskOut_1_0_7(dataModule_io_maskOut_1_0_7),
    .io_maskOut_1_1_0(dataModule_io_maskOut_1_1_0),
    .io_maskOut_1_1_1(dataModule_io_maskOut_1_1_1),
    .io_maskOut_1_1_2(dataModule_io_maskOut_1_1_2),
    .io_maskOut_1_1_3(dataModule_io_maskOut_1_1_3),
    .io_maskOut_1_1_4(dataModule_io_maskOut_1_1_4),
    .io_maskOut_1_1_5(dataModule_io_maskOut_1_1_5),
    .io_maskOut_1_1_6(dataModule_io_maskOut_1_1_6),
    .io_maskOut_1_1_7(dataModule_io_maskOut_1_1_7),
    .io_maskOut_1_2_0(dataModule_io_maskOut_1_2_0),
    .io_maskOut_1_2_1(dataModule_io_maskOut_1_2_1),
    .io_maskOut_1_2_2(dataModule_io_maskOut_1_2_2),
    .io_maskOut_1_2_3(dataModule_io_maskOut_1_2_3),
    .io_maskOut_1_2_4(dataModule_io_maskOut_1_2_4),
    .io_maskOut_1_2_5(dataModule_io_maskOut_1_2_5),
    .io_maskOut_1_2_6(dataModule_io_maskOut_1_2_6),
    .io_maskOut_1_2_7(dataModule_io_maskOut_1_2_7),
    .io_maskOut_1_3_0(dataModule_io_maskOut_1_3_0),
    .io_maskOut_1_3_1(dataModule_io_maskOut_1_3_1),
    .io_maskOut_1_3_2(dataModule_io_maskOut_1_3_2),
    .io_maskOut_1_3_3(dataModule_io_maskOut_1_3_3),
    .io_maskOut_1_3_4(dataModule_io_maskOut_1_3_4),
    .io_maskOut_1_3_5(dataModule_io_maskOut_1_3_5),
    .io_maskOut_1_3_6(dataModule_io_maskOut_1_3_6),
    .io_maskOut_1_3_7(dataModule_io_maskOut_1_3_7),
    .io_maskOut_1_4_0(dataModule_io_maskOut_1_4_0),
    .io_maskOut_1_4_1(dataModule_io_maskOut_1_4_1),
    .io_maskOut_1_4_2(dataModule_io_maskOut_1_4_2),
    .io_maskOut_1_4_3(dataModule_io_maskOut_1_4_3),
    .io_maskOut_1_4_4(dataModule_io_maskOut_1_4_4),
    .io_maskOut_1_4_5(dataModule_io_maskOut_1_4_5),
    .io_maskOut_1_4_6(dataModule_io_maskOut_1_4_6),
    .io_maskOut_1_4_7(dataModule_io_maskOut_1_4_7),
    .io_maskOut_1_5_0(dataModule_io_maskOut_1_5_0),
    .io_maskOut_1_5_1(dataModule_io_maskOut_1_5_1),
    .io_maskOut_1_5_2(dataModule_io_maskOut_1_5_2),
    .io_maskOut_1_5_3(dataModule_io_maskOut_1_5_3),
    .io_maskOut_1_5_4(dataModule_io_maskOut_1_5_4),
    .io_maskOut_1_5_5(dataModule_io_maskOut_1_5_5),
    .io_maskOut_1_5_6(dataModule_io_maskOut_1_5_6),
    .io_maskOut_1_5_7(dataModule_io_maskOut_1_5_7),
    .io_maskOut_1_6_0(dataModule_io_maskOut_1_6_0),
    .io_maskOut_1_6_1(dataModule_io_maskOut_1_6_1),
    .io_maskOut_1_6_2(dataModule_io_maskOut_1_6_2),
    .io_maskOut_1_6_3(dataModule_io_maskOut_1_6_3),
    .io_maskOut_1_6_4(dataModule_io_maskOut_1_6_4),
    .io_maskOut_1_6_5(dataModule_io_maskOut_1_6_5),
    .io_maskOut_1_6_6(dataModule_io_maskOut_1_6_6),
    .io_maskOut_1_6_7(dataModule_io_maskOut_1_6_7),
    .io_maskOut_1_7_0(dataModule_io_maskOut_1_7_0),
    .io_maskOut_1_7_1(dataModule_io_maskOut_1_7_1),
    .io_maskOut_1_7_2(dataModule_io_maskOut_1_7_2),
    .io_maskOut_1_7_3(dataModule_io_maskOut_1_7_3),
    .io_maskOut_1_7_4(dataModule_io_maskOut_1_7_4),
    .io_maskOut_1_7_5(dataModule_io_maskOut_1_7_5),
    .io_maskOut_1_7_6(dataModule_io_maskOut_1_7_6),
    .io_maskOut_1_7_7(dataModule_io_maskOut_1_7_7),
    .io_maskOut_2_0_0(dataModule_io_maskOut_2_0_0),
    .io_maskOut_2_0_1(dataModule_io_maskOut_2_0_1),
    .io_maskOut_2_0_2(dataModule_io_maskOut_2_0_2),
    .io_maskOut_2_0_3(dataModule_io_maskOut_2_0_3),
    .io_maskOut_2_0_4(dataModule_io_maskOut_2_0_4),
    .io_maskOut_2_0_5(dataModule_io_maskOut_2_0_5),
    .io_maskOut_2_0_6(dataModule_io_maskOut_2_0_6),
    .io_maskOut_2_0_7(dataModule_io_maskOut_2_0_7),
    .io_maskOut_2_1_0(dataModule_io_maskOut_2_1_0),
    .io_maskOut_2_1_1(dataModule_io_maskOut_2_1_1),
    .io_maskOut_2_1_2(dataModule_io_maskOut_2_1_2),
    .io_maskOut_2_1_3(dataModule_io_maskOut_2_1_3),
    .io_maskOut_2_1_4(dataModule_io_maskOut_2_1_4),
    .io_maskOut_2_1_5(dataModule_io_maskOut_2_1_5),
    .io_maskOut_2_1_6(dataModule_io_maskOut_2_1_6),
    .io_maskOut_2_1_7(dataModule_io_maskOut_2_1_7),
    .io_maskOut_2_2_0(dataModule_io_maskOut_2_2_0),
    .io_maskOut_2_2_1(dataModule_io_maskOut_2_2_1),
    .io_maskOut_2_2_2(dataModule_io_maskOut_2_2_2),
    .io_maskOut_2_2_3(dataModule_io_maskOut_2_2_3),
    .io_maskOut_2_2_4(dataModule_io_maskOut_2_2_4),
    .io_maskOut_2_2_5(dataModule_io_maskOut_2_2_5),
    .io_maskOut_2_2_6(dataModule_io_maskOut_2_2_6),
    .io_maskOut_2_2_7(dataModule_io_maskOut_2_2_7),
    .io_maskOut_2_3_0(dataModule_io_maskOut_2_3_0),
    .io_maskOut_2_3_1(dataModule_io_maskOut_2_3_1),
    .io_maskOut_2_3_2(dataModule_io_maskOut_2_3_2),
    .io_maskOut_2_3_3(dataModule_io_maskOut_2_3_3),
    .io_maskOut_2_3_4(dataModule_io_maskOut_2_3_4),
    .io_maskOut_2_3_5(dataModule_io_maskOut_2_3_5),
    .io_maskOut_2_3_6(dataModule_io_maskOut_2_3_6),
    .io_maskOut_2_3_7(dataModule_io_maskOut_2_3_7),
    .io_maskOut_2_4_0(dataModule_io_maskOut_2_4_0),
    .io_maskOut_2_4_1(dataModule_io_maskOut_2_4_1),
    .io_maskOut_2_4_2(dataModule_io_maskOut_2_4_2),
    .io_maskOut_2_4_3(dataModule_io_maskOut_2_4_3),
    .io_maskOut_2_4_4(dataModule_io_maskOut_2_4_4),
    .io_maskOut_2_4_5(dataModule_io_maskOut_2_4_5),
    .io_maskOut_2_4_6(dataModule_io_maskOut_2_4_6),
    .io_maskOut_2_4_7(dataModule_io_maskOut_2_4_7),
    .io_maskOut_2_5_0(dataModule_io_maskOut_2_5_0),
    .io_maskOut_2_5_1(dataModule_io_maskOut_2_5_1),
    .io_maskOut_2_5_2(dataModule_io_maskOut_2_5_2),
    .io_maskOut_2_5_3(dataModule_io_maskOut_2_5_3),
    .io_maskOut_2_5_4(dataModule_io_maskOut_2_5_4),
    .io_maskOut_2_5_5(dataModule_io_maskOut_2_5_5),
    .io_maskOut_2_5_6(dataModule_io_maskOut_2_5_6),
    .io_maskOut_2_5_7(dataModule_io_maskOut_2_5_7),
    .io_maskOut_2_6_0(dataModule_io_maskOut_2_6_0),
    .io_maskOut_2_6_1(dataModule_io_maskOut_2_6_1),
    .io_maskOut_2_6_2(dataModule_io_maskOut_2_6_2),
    .io_maskOut_2_6_3(dataModule_io_maskOut_2_6_3),
    .io_maskOut_2_6_4(dataModule_io_maskOut_2_6_4),
    .io_maskOut_2_6_5(dataModule_io_maskOut_2_6_5),
    .io_maskOut_2_6_6(dataModule_io_maskOut_2_6_6),
    .io_maskOut_2_6_7(dataModule_io_maskOut_2_6_7),
    .io_maskOut_2_7_0(dataModule_io_maskOut_2_7_0),
    .io_maskOut_2_7_1(dataModule_io_maskOut_2_7_1),
    .io_maskOut_2_7_2(dataModule_io_maskOut_2_7_2),
    .io_maskOut_2_7_3(dataModule_io_maskOut_2_7_3),
    .io_maskOut_2_7_4(dataModule_io_maskOut_2_7_4),
    .io_maskOut_2_7_5(dataModule_io_maskOut_2_7_5),
    .io_maskOut_2_7_6(dataModule_io_maskOut_2_7_6),
    .io_maskOut_2_7_7(dataModule_io_maskOut_2_7_7),
    .io_maskOut_3_0_0(dataModule_io_maskOut_3_0_0),
    .io_maskOut_3_0_1(dataModule_io_maskOut_3_0_1),
    .io_maskOut_3_0_2(dataModule_io_maskOut_3_0_2),
    .io_maskOut_3_0_3(dataModule_io_maskOut_3_0_3),
    .io_maskOut_3_0_4(dataModule_io_maskOut_3_0_4),
    .io_maskOut_3_0_5(dataModule_io_maskOut_3_0_5),
    .io_maskOut_3_0_6(dataModule_io_maskOut_3_0_6),
    .io_maskOut_3_0_7(dataModule_io_maskOut_3_0_7),
    .io_maskOut_3_1_0(dataModule_io_maskOut_3_1_0),
    .io_maskOut_3_1_1(dataModule_io_maskOut_3_1_1),
    .io_maskOut_3_1_2(dataModule_io_maskOut_3_1_2),
    .io_maskOut_3_1_3(dataModule_io_maskOut_3_1_3),
    .io_maskOut_3_1_4(dataModule_io_maskOut_3_1_4),
    .io_maskOut_3_1_5(dataModule_io_maskOut_3_1_5),
    .io_maskOut_3_1_6(dataModule_io_maskOut_3_1_6),
    .io_maskOut_3_1_7(dataModule_io_maskOut_3_1_7),
    .io_maskOut_3_2_0(dataModule_io_maskOut_3_2_0),
    .io_maskOut_3_2_1(dataModule_io_maskOut_3_2_1),
    .io_maskOut_3_2_2(dataModule_io_maskOut_3_2_2),
    .io_maskOut_3_2_3(dataModule_io_maskOut_3_2_3),
    .io_maskOut_3_2_4(dataModule_io_maskOut_3_2_4),
    .io_maskOut_3_2_5(dataModule_io_maskOut_3_2_5),
    .io_maskOut_3_2_6(dataModule_io_maskOut_3_2_6),
    .io_maskOut_3_2_7(dataModule_io_maskOut_3_2_7),
    .io_maskOut_3_3_0(dataModule_io_maskOut_3_3_0),
    .io_maskOut_3_3_1(dataModule_io_maskOut_3_3_1),
    .io_maskOut_3_3_2(dataModule_io_maskOut_3_3_2),
    .io_maskOut_3_3_3(dataModule_io_maskOut_3_3_3),
    .io_maskOut_3_3_4(dataModule_io_maskOut_3_3_4),
    .io_maskOut_3_3_5(dataModule_io_maskOut_3_3_5),
    .io_maskOut_3_3_6(dataModule_io_maskOut_3_3_6),
    .io_maskOut_3_3_7(dataModule_io_maskOut_3_3_7),
    .io_maskOut_3_4_0(dataModule_io_maskOut_3_4_0),
    .io_maskOut_3_4_1(dataModule_io_maskOut_3_4_1),
    .io_maskOut_3_4_2(dataModule_io_maskOut_3_4_2),
    .io_maskOut_3_4_3(dataModule_io_maskOut_3_4_3),
    .io_maskOut_3_4_4(dataModule_io_maskOut_3_4_4),
    .io_maskOut_3_4_5(dataModule_io_maskOut_3_4_5),
    .io_maskOut_3_4_6(dataModule_io_maskOut_3_4_6),
    .io_maskOut_3_4_7(dataModule_io_maskOut_3_4_7),
    .io_maskOut_3_5_0(dataModule_io_maskOut_3_5_0),
    .io_maskOut_3_5_1(dataModule_io_maskOut_3_5_1),
    .io_maskOut_3_5_2(dataModule_io_maskOut_3_5_2),
    .io_maskOut_3_5_3(dataModule_io_maskOut_3_5_3),
    .io_maskOut_3_5_4(dataModule_io_maskOut_3_5_4),
    .io_maskOut_3_5_5(dataModule_io_maskOut_3_5_5),
    .io_maskOut_3_5_6(dataModule_io_maskOut_3_5_6),
    .io_maskOut_3_5_7(dataModule_io_maskOut_3_5_7),
    .io_maskOut_3_6_0(dataModule_io_maskOut_3_6_0),
    .io_maskOut_3_6_1(dataModule_io_maskOut_3_6_1),
    .io_maskOut_3_6_2(dataModule_io_maskOut_3_6_2),
    .io_maskOut_3_6_3(dataModule_io_maskOut_3_6_3),
    .io_maskOut_3_6_4(dataModule_io_maskOut_3_6_4),
    .io_maskOut_3_6_5(dataModule_io_maskOut_3_6_5),
    .io_maskOut_3_6_6(dataModule_io_maskOut_3_6_6),
    .io_maskOut_3_6_7(dataModule_io_maskOut_3_6_7),
    .io_maskOut_3_7_0(dataModule_io_maskOut_3_7_0),
    .io_maskOut_3_7_1(dataModule_io_maskOut_3_7_1),
    .io_maskOut_3_7_2(dataModule_io_maskOut_3_7_2),
    .io_maskOut_3_7_3(dataModule_io_maskOut_3_7_3),
    .io_maskOut_3_7_4(dataModule_io_maskOut_3_7_4),
    .io_maskOut_3_7_5(dataModule_io_maskOut_3_7_5),
    .io_maskOut_3_7_6(dataModule_io_maskOut_3_7_6),
    .io_maskOut_3_7_7(dataModule_io_maskOut_3_7_7),
    .io_maskOut_4_0_0(dataModule_io_maskOut_4_0_0),
    .io_maskOut_4_0_1(dataModule_io_maskOut_4_0_1),
    .io_maskOut_4_0_2(dataModule_io_maskOut_4_0_2),
    .io_maskOut_4_0_3(dataModule_io_maskOut_4_0_3),
    .io_maskOut_4_0_4(dataModule_io_maskOut_4_0_4),
    .io_maskOut_4_0_5(dataModule_io_maskOut_4_0_5),
    .io_maskOut_4_0_6(dataModule_io_maskOut_4_0_6),
    .io_maskOut_4_0_7(dataModule_io_maskOut_4_0_7),
    .io_maskOut_4_1_0(dataModule_io_maskOut_4_1_0),
    .io_maskOut_4_1_1(dataModule_io_maskOut_4_1_1),
    .io_maskOut_4_1_2(dataModule_io_maskOut_4_1_2),
    .io_maskOut_4_1_3(dataModule_io_maskOut_4_1_3),
    .io_maskOut_4_1_4(dataModule_io_maskOut_4_1_4),
    .io_maskOut_4_1_5(dataModule_io_maskOut_4_1_5),
    .io_maskOut_4_1_6(dataModule_io_maskOut_4_1_6),
    .io_maskOut_4_1_7(dataModule_io_maskOut_4_1_7),
    .io_maskOut_4_2_0(dataModule_io_maskOut_4_2_0),
    .io_maskOut_4_2_1(dataModule_io_maskOut_4_2_1),
    .io_maskOut_4_2_2(dataModule_io_maskOut_4_2_2),
    .io_maskOut_4_2_3(dataModule_io_maskOut_4_2_3),
    .io_maskOut_4_2_4(dataModule_io_maskOut_4_2_4),
    .io_maskOut_4_2_5(dataModule_io_maskOut_4_2_5),
    .io_maskOut_4_2_6(dataModule_io_maskOut_4_2_6),
    .io_maskOut_4_2_7(dataModule_io_maskOut_4_2_7),
    .io_maskOut_4_3_0(dataModule_io_maskOut_4_3_0),
    .io_maskOut_4_3_1(dataModule_io_maskOut_4_3_1),
    .io_maskOut_4_3_2(dataModule_io_maskOut_4_3_2),
    .io_maskOut_4_3_3(dataModule_io_maskOut_4_3_3),
    .io_maskOut_4_3_4(dataModule_io_maskOut_4_3_4),
    .io_maskOut_4_3_5(dataModule_io_maskOut_4_3_5),
    .io_maskOut_4_3_6(dataModule_io_maskOut_4_3_6),
    .io_maskOut_4_3_7(dataModule_io_maskOut_4_3_7),
    .io_maskOut_4_4_0(dataModule_io_maskOut_4_4_0),
    .io_maskOut_4_4_1(dataModule_io_maskOut_4_4_1),
    .io_maskOut_4_4_2(dataModule_io_maskOut_4_4_2),
    .io_maskOut_4_4_3(dataModule_io_maskOut_4_4_3),
    .io_maskOut_4_4_4(dataModule_io_maskOut_4_4_4),
    .io_maskOut_4_4_5(dataModule_io_maskOut_4_4_5),
    .io_maskOut_4_4_6(dataModule_io_maskOut_4_4_6),
    .io_maskOut_4_4_7(dataModule_io_maskOut_4_4_7),
    .io_maskOut_4_5_0(dataModule_io_maskOut_4_5_0),
    .io_maskOut_4_5_1(dataModule_io_maskOut_4_5_1),
    .io_maskOut_4_5_2(dataModule_io_maskOut_4_5_2),
    .io_maskOut_4_5_3(dataModule_io_maskOut_4_5_3),
    .io_maskOut_4_5_4(dataModule_io_maskOut_4_5_4),
    .io_maskOut_4_5_5(dataModule_io_maskOut_4_5_5),
    .io_maskOut_4_5_6(dataModule_io_maskOut_4_5_6),
    .io_maskOut_4_5_7(dataModule_io_maskOut_4_5_7),
    .io_maskOut_4_6_0(dataModule_io_maskOut_4_6_0),
    .io_maskOut_4_6_1(dataModule_io_maskOut_4_6_1),
    .io_maskOut_4_6_2(dataModule_io_maskOut_4_6_2),
    .io_maskOut_4_6_3(dataModule_io_maskOut_4_6_3),
    .io_maskOut_4_6_4(dataModule_io_maskOut_4_6_4),
    .io_maskOut_4_6_5(dataModule_io_maskOut_4_6_5),
    .io_maskOut_4_6_6(dataModule_io_maskOut_4_6_6),
    .io_maskOut_4_6_7(dataModule_io_maskOut_4_6_7),
    .io_maskOut_4_7_0(dataModule_io_maskOut_4_7_0),
    .io_maskOut_4_7_1(dataModule_io_maskOut_4_7_1),
    .io_maskOut_4_7_2(dataModule_io_maskOut_4_7_2),
    .io_maskOut_4_7_3(dataModule_io_maskOut_4_7_3),
    .io_maskOut_4_7_4(dataModule_io_maskOut_4_7_4),
    .io_maskOut_4_7_5(dataModule_io_maskOut_4_7_5),
    .io_maskOut_4_7_6(dataModule_io_maskOut_4_7_6),
    .io_maskOut_4_7_7(dataModule_io_maskOut_4_7_7),
    .io_maskOut_5_0_0(dataModule_io_maskOut_5_0_0),
    .io_maskOut_5_0_1(dataModule_io_maskOut_5_0_1),
    .io_maskOut_5_0_2(dataModule_io_maskOut_5_0_2),
    .io_maskOut_5_0_3(dataModule_io_maskOut_5_0_3),
    .io_maskOut_5_0_4(dataModule_io_maskOut_5_0_4),
    .io_maskOut_5_0_5(dataModule_io_maskOut_5_0_5),
    .io_maskOut_5_0_6(dataModule_io_maskOut_5_0_6),
    .io_maskOut_5_0_7(dataModule_io_maskOut_5_0_7),
    .io_maskOut_5_1_0(dataModule_io_maskOut_5_1_0),
    .io_maskOut_5_1_1(dataModule_io_maskOut_5_1_1),
    .io_maskOut_5_1_2(dataModule_io_maskOut_5_1_2),
    .io_maskOut_5_1_3(dataModule_io_maskOut_5_1_3),
    .io_maskOut_5_1_4(dataModule_io_maskOut_5_1_4),
    .io_maskOut_5_1_5(dataModule_io_maskOut_5_1_5),
    .io_maskOut_5_1_6(dataModule_io_maskOut_5_1_6),
    .io_maskOut_5_1_7(dataModule_io_maskOut_5_1_7),
    .io_maskOut_5_2_0(dataModule_io_maskOut_5_2_0),
    .io_maskOut_5_2_1(dataModule_io_maskOut_5_2_1),
    .io_maskOut_5_2_2(dataModule_io_maskOut_5_2_2),
    .io_maskOut_5_2_3(dataModule_io_maskOut_5_2_3),
    .io_maskOut_5_2_4(dataModule_io_maskOut_5_2_4),
    .io_maskOut_5_2_5(dataModule_io_maskOut_5_2_5),
    .io_maskOut_5_2_6(dataModule_io_maskOut_5_2_6),
    .io_maskOut_5_2_7(dataModule_io_maskOut_5_2_7),
    .io_maskOut_5_3_0(dataModule_io_maskOut_5_3_0),
    .io_maskOut_5_3_1(dataModule_io_maskOut_5_3_1),
    .io_maskOut_5_3_2(dataModule_io_maskOut_5_3_2),
    .io_maskOut_5_3_3(dataModule_io_maskOut_5_3_3),
    .io_maskOut_5_3_4(dataModule_io_maskOut_5_3_4),
    .io_maskOut_5_3_5(dataModule_io_maskOut_5_3_5),
    .io_maskOut_5_3_6(dataModule_io_maskOut_5_3_6),
    .io_maskOut_5_3_7(dataModule_io_maskOut_5_3_7),
    .io_maskOut_5_4_0(dataModule_io_maskOut_5_4_0),
    .io_maskOut_5_4_1(dataModule_io_maskOut_5_4_1),
    .io_maskOut_5_4_2(dataModule_io_maskOut_5_4_2),
    .io_maskOut_5_4_3(dataModule_io_maskOut_5_4_3),
    .io_maskOut_5_4_4(dataModule_io_maskOut_5_4_4),
    .io_maskOut_5_4_5(dataModule_io_maskOut_5_4_5),
    .io_maskOut_5_4_6(dataModule_io_maskOut_5_4_6),
    .io_maskOut_5_4_7(dataModule_io_maskOut_5_4_7),
    .io_maskOut_5_5_0(dataModule_io_maskOut_5_5_0),
    .io_maskOut_5_5_1(dataModule_io_maskOut_5_5_1),
    .io_maskOut_5_5_2(dataModule_io_maskOut_5_5_2),
    .io_maskOut_5_5_3(dataModule_io_maskOut_5_5_3),
    .io_maskOut_5_5_4(dataModule_io_maskOut_5_5_4),
    .io_maskOut_5_5_5(dataModule_io_maskOut_5_5_5),
    .io_maskOut_5_5_6(dataModule_io_maskOut_5_5_6),
    .io_maskOut_5_5_7(dataModule_io_maskOut_5_5_7),
    .io_maskOut_5_6_0(dataModule_io_maskOut_5_6_0),
    .io_maskOut_5_6_1(dataModule_io_maskOut_5_6_1),
    .io_maskOut_5_6_2(dataModule_io_maskOut_5_6_2),
    .io_maskOut_5_6_3(dataModule_io_maskOut_5_6_3),
    .io_maskOut_5_6_4(dataModule_io_maskOut_5_6_4),
    .io_maskOut_5_6_5(dataModule_io_maskOut_5_6_5),
    .io_maskOut_5_6_6(dataModule_io_maskOut_5_6_6),
    .io_maskOut_5_6_7(dataModule_io_maskOut_5_6_7),
    .io_maskOut_5_7_0(dataModule_io_maskOut_5_7_0),
    .io_maskOut_5_7_1(dataModule_io_maskOut_5_7_1),
    .io_maskOut_5_7_2(dataModule_io_maskOut_5_7_2),
    .io_maskOut_5_7_3(dataModule_io_maskOut_5_7_3),
    .io_maskOut_5_7_4(dataModule_io_maskOut_5_7_4),
    .io_maskOut_5_7_5(dataModule_io_maskOut_5_7_5),
    .io_maskOut_5_7_6(dataModule_io_maskOut_5_7_6),
    .io_maskOut_5_7_7(dataModule_io_maskOut_5_7_7),
    .io_maskOut_6_0_0(dataModule_io_maskOut_6_0_0),
    .io_maskOut_6_0_1(dataModule_io_maskOut_6_0_1),
    .io_maskOut_6_0_2(dataModule_io_maskOut_6_0_2),
    .io_maskOut_6_0_3(dataModule_io_maskOut_6_0_3),
    .io_maskOut_6_0_4(dataModule_io_maskOut_6_0_4),
    .io_maskOut_6_0_5(dataModule_io_maskOut_6_0_5),
    .io_maskOut_6_0_6(dataModule_io_maskOut_6_0_6),
    .io_maskOut_6_0_7(dataModule_io_maskOut_6_0_7),
    .io_maskOut_6_1_0(dataModule_io_maskOut_6_1_0),
    .io_maskOut_6_1_1(dataModule_io_maskOut_6_1_1),
    .io_maskOut_6_1_2(dataModule_io_maskOut_6_1_2),
    .io_maskOut_6_1_3(dataModule_io_maskOut_6_1_3),
    .io_maskOut_6_1_4(dataModule_io_maskOut_6_1_4),
    .io_maskOut_6_1_5(dataModule_io_maskOut_6_1_5),
    .io_maskOut_6_1_6(dataModule_io_maskOut_6_1_6),
    .io_maskOut_6_1_7(dataModule_io_maskOut_6_1_7),
    .io_maskOut_6_2_0(dataModule_io_maskOut_6_2_0),
    .io_maskOut_6_2_1(dataModule_io_maskOut_6_2_1),
    .io_maskOut_6_2_2(dataModule_io_maskOut_6_2_2),
    .io_maskOut_6_2_3(dataModule_io_maskOut_6_2_3),
    .io_maskOut_6_2_4(dataModule_io_maskOut_6_2_4),
    .io_maskOut_6_2_5(dataModule_io_maskOut_6_2_5),
    .io_maskOut_6_2_6(dataModule_io_maskOut_6_2_6),
    .io_maskOut_6_2_7(dataModule_io_maskOut_6_2_7),
    .io_maskOut_6_3_0(dataModule_io_maskOut_6_3_0),
    .io_maskOut_6_3_1(dataModule_io_maskOut_6_3_1),
    .io_maskOut_6_3_2(dataModule_io_maskOut_6_3_2),
    .io_maskOut_6_3_3(dataModule_io_maskOut_6_3_3),
    .io_maskOut_6_3_4(dataModule_io_maskOut_6_3_4),
    .io_maskOut_6_3_5(dataModule_io_maskOut_6_3_5),
    .io_maskOut_6_3_6(dataModule_io_maskOut_6_3_6),
    .io_maskOut_6_3_7(dataModule_io_maskOut_6_3_7),
    .io_maskOut_6_4_0(dataModule_io_maskOut_6_4_0),
    .io_maskOut_6_4_1(dataModule_io_maskOut_6_4_1),
    .io_maskOut_6_4_2(dataModule_io_maskOut_6_4_2),
    .io_maskOut_6_4_3(dataModule_io_maskOut_6_4_3),
    .io_maskOut_6_4_4(dataModule_io_maskOut_6_4_4),
    .io_maskOut_6_4_5(dataModule_io_maskOut_6_4_5),
    .io_maskOut_6_4_6(dataModule_io_maskOut_6_4_6),
    .io_maskOut_6_4_7(dataModule_io_maskOut_6_4_7),
    .io_maskOut_6_5_0(dataModule_io_maskOut_6_5_0),
    .io_maskOut_6_5_1(dataModule_io_maskOut_6_5_1),
    .io_maskOut_6_5_2(dataModule_io_maskOut_6_5_2),
    .io_maskOut_6_5_3(dataModule_io_maskOut_6_5_3),
    .io_maskOut_6_5_4(dataModule_io_maskOut_6_5_4),
    .io_maskOut_6_5_5(dataModule_io_maskOut_6_5_5),
    .io_maskOut_6_5_6(dataModule_io_maskOut_6_5_6),
    .io_maskOut_6_5_7(dataModule_io_maskOut_6_5_7),
    .io_maskOut_6_6_0(dataModule_io_maskOut_6_6_0),
    .io_maskOut_6_6_1(dataModule_io_maskOut_6_6_1),
    .io_maskOut_6_6_2(dataModule_io_maskOut_6_6_2),
    .io_maskOut_6_6_3(dataModule_io_maskOut_6_6_3),
    .io_maskOut_6_6_4(dataModule_io_maskOut_6_6_4),
    .io_maskOut_6_6_5(dataModule_io_maskOut_6_6_5),
    .io_maskOut_6_6_6(dataModule_io_maskOut_6_6_6),
    .io_maskOut_6_6_7(dataModule_io_maskOut_6_6_7),
    .io_maskOut_6_7_0(dataModule_io_maskOut_6_7_0),
    .io_maskOut_6_7_1(dataModule_io_maskOut_6_7_1),
    .io_maskOut_6_7_2(dataModule_io_maskOut_6_7_2),
    .io_maskOut_6_7_3(dataModule_io_maskOut_6_7_3),
    .io_maskOut_6_7_4(dataModule_io_maskOut_6_7_4),
    .io_maskOut_6_7_5(dataModule_io_maskOut_6_7_5),
    .io_maskOut_6_7_6(dataModule_io_maskOut_6_7_6),
    .io_maskOut_6_7_7(dataModule_io_maskOut_6_7_7),
    .io_maskOut_7_0_0(dataModule_io_maskOut_7_0_0),
    .io_maskOut_7_0_1(dataModule_io_maskOut_7_0_1),
    .io_maskOut_7_0_2(dataModule_io_maskOut_7_0_2),
    .io_maskOut_7_0_3(dataModule_io_maskOut_7_0_3),
    .io_maskOut_7_0_4(dataModule_io_maskOut_7_0_4),
    .io_maskOut_7_0_5(dataModule_io_maskOut_7_0_5),
    .io_maskOut_7_0_6(dataModule_io_maskOut_7_0_6),
    .io_maskOut_7_0_7(dataModule_io_maskOut_7_0_7),
    .io_maskOut_7_1_0(dataModule_io_maskOut_7_1_0),
    .io_maskOut_7_1_1(dataModule_io_maskOut_7_1_1),
    .io_maskOut_7_1_2(dataModule_io_maskOut_7_1_2),
    .io_maskOut_7_1_3(dataModule_io_maskOut_7_1_3),
    .io_maskOut_7_1_4(dataModule_io_maskOut_7_1_4),
    .io_maskOut_7_1_5(dataModule_io_maskOut_7_1_5),
    .io_maskOut_7_1_6(dataModule_io_maskOut_7_1_6),
    .io_maskOut_7_1_7(dataModule_io_maskOut_7_1_7),
    .io_maskOut_7_2_0(dataModule_io_maskOut_7_2_0),
    .io_maskOut_7_2_1(dataModule_io_maskOut_7_2_1),
    .io_maskOut_7_2_2(dataModule_io_maskOut_7_2_2),
    .io_maskOut_7_2_3(dataModule_io_maskOut_7_2_3),
    .io_maskOut_7_2_4(dataModule_io_maskOut_7_2_4),
    .io_maskOut_7_2_5(dataModule_io_maskOut_7_2_5),
    .io_maskOut_7_2_6(dataModule_io_maskOut_7_2_6),
    .io_maskOut_7_2_7(dataModule_io_maskOut_7_2_7),
    .io_maskOut_7_3_0(dataModule_io_maskOut_7_3_0),
    .io_maskOut_7_3_1(dataModule_io_maskOut_7_3_1),
    .io_maskOut_7_3_2(dataModule_io_maskOut_7_3_2),
    .io_maskOut_7_3_3(dataModule_io_maskOut_7_3_3),
    .io_maskOut_7_3_4(dataModule_io_maskOut_7_3_4),
    .io_maskOut_7_3_5(dataModule_io_maskOut_7_3_5),
    .io_maskOut_7_3_6(dataModule_io_maskOut_7_3_6),
    .io_maskOut_7_3_7(dataModule_io_maskOut_7_3_7),
    .io_maskOut_7_4_0(dataModule_io_maskOut_7_4_0),
    .io_maskOut_7_4_1(dataModule_io_maskOut_7_4_1),
    .io_maskOut_7_4_2(dataModule_io_maskOut_7_4_2),
    .io_maskOut_7_4_3(dataModule_io_maskOut_7_4_3),
    .io_maskOut_7_4_4(dataModule_io_maskOut_7_4_4),
    .io_maskOut_7_4_5(dataModule_io_maskOut_7_4_5),
    .io_maskOut_7_4_6(dataModule_io_maskOut_7_4_6),
    .io_maskOut_7_4_7(dataModule_io_maskOut_7_4_7),
    .io_maskOut_7_5_0(dataModule_io_maskOut_7_5_0),
    .io_maskOut_7_5_1(dataModule_io_maskOut_7_5_1),
    .io_maskOut_7_5_2(dataModule_io_maskOut_7_5_2),
    .io_maskOut_7_5_3(dataModule_io_maskOut_7_5_3),
    .io_maskOut_7_5_4(dataModule_io_maskOut_7_5_4),
    .io_maskOut_7_5_5(dataModule_io_maskOut_7_5_5),
    .io_maskOut_7_5_6(dataModule_io_maskOut_7_5_6),
    .io_maskOut_7_5_7(dataModule_io_maskOut_7_5_7),
    .io_maskOut_7_6_0(dataModule_io_maskOut_7_6_0),
    .io_maskOut_7_6_1(dataModule_io_maskOut_7_6_1),
    .io_maskOut_7_6_2(dataModule_io_maskOut_7_6_2),
    .io_maskOut_7_6_3(dataModule_io_maskOut_7_6_3),
    .io_maskOut_7_6_4(dataModule_io_maskOut_7_6_4),
    .io_maskOut_7_6_5(dataModule_io_maskOut_7_6_5),
    .io_maskOut_7_6_6(dataModule_io_maskOut_7_6_6),
    .io_maskOut_7_6_7(dataModule_io_maskOut_7_6_7),
    .io_maskOut_7_7_0(dataModule_io_maskOut_7_7_0),
    .io_maskOut_7_7_1(dataModule_io_maskOut_7_7_1),
    .io_maskOut_7_7_2(dataModule_io_maskOut_7_7_2),
    .io_maskOut_7_7_3(dataModule_io_maskOut_7_7_3),
    .io_maskOut_7_7_4(dataModule_io_maskOut_7_7_4),
    .io_maskOut_7_7_5(dataModule_io_maskOut_7_7_5),
    .io_maskOut_7_7_6(dataModule_io_maskOut_7_7_6),
    .io_maskOut_7_7_7(dataModule_io_maskOut_7_7_7),
    .io_maskOut_8_0_0(dataModule_io_maskOut_8_0_0),
    .io_maskOut_8_0_1(dataModule_io_maskOut_8_0_1),
    .io_maskOut_8_0_2(dataModule_io_maskOut_8_0_2),
    .io_maskOut_8_0_3(dataModule_io_maskOut_8_0_3),
    .io_maskOut_8_0_4(dataModule_io_maskOut_8_0_4),
    .io_maskOut_8_0_5(dataModule_io_maskOut_8_0_5),
    .io_maskOut_8_0_6(dataModule_io_maskOut_8_0_6),
    .io_maskOut_8_0_7(dataModule_io_maskOut_8_0_7),
    .io_maskOut_8_1_0(dataModule_io_maskOut_8_1_0),
    .io_maskOut_8_1_1(dataModule_io_maskOut_8_1_1),
    .io_maskOut_8_1_2(dataModule_io_maskOut_8_1_2),
    .io_maskOut_8_1_3(dataModule_io_maskOut_8_1_3),
    .io_maskOut_8_1_4(dataModule_io_maskOut_8_1_4),
    .io_maskOut_8_1_5(dataModule_io_maskOut_8_1_5),
    .io_maskOut_8_1_6(dataModule_io_maskOut_8_1_6),
    .io_maskOut_8_1_7(dataModule_io_maskOut_8_1_7),
    .io_maskOut_8_2_0(dataModule_io_maskOut_8_2_0),
    .io_maskOut_8_2_1(dataModule_io_maskOut_8_2_1),
    .io_maskOut_8_2_2(dataModule_io_maskOut_8_2_2),
    .io_maskOut_8_2_3(dataModule_io_maskOut_8_2_3),
    .io_maskOut_8_2_4(dataModule_io_maskOut_8_2_4),
    .io_maskOut_8_2_5(dataModule_io_maskOut_8_2_5),
    .io_maskOut_8_2_6(dataModule_io_maskOut_8_2_6),
    .io_maskOut_8_2_7(dataModule_io_maskOut_8_2_7),
    .io_maskOut_8_3_0(dataModule_io_maskOut_8_3_0),
    .io_maskOut_8_3_1(dataModule_io_maskOut_8_3_1),
    .io_maskOut_8_3_2(dataModule_io_maskOut_8_3_2),
    .io_maskOut_8_3_3(dataModule_io_maskOut_8_3_3),
    .io_maskOut_8_3_4(dataModule_io_maskOut_8_3_4),
    .io_maskOut_8_3_5(dataModule_io_maskOut_8_3_5),
    .io_maskOut_8_3_6(dataModule_io_maskOut_8_3_6),
    .io_maskOut_8_3_7(dataModule_io_maskOut_8_3_7),
    .io_maskOut_8_4_0(dataModule_io_maskOut_8_4_0),
    .io_maskOut_8_4_1(dataModule_io_maskOut_8_4_1),
    .io_maskOut_8_4_2(dataModule_io_maskOut_8_4_2),
    .io_maskOut_8_4_3(dataModule_io_maskOut_8_4_3),
    .io_maskOut_8_4_4(dataModule_io_maskOut_8_4_4),
    .io_maskOut_8_4_5(dataModule_io_maskOut_8_4_5),
    .io_maskOut_8_4_6(dataModule_io_maskOut_8_4_6),
    .io_maskOut_8_4_7(dataModule_io_maskOut_8_4_7),
    .io_maskOut_8_5_0(dataModule_io_maskOut_8_5_0),
    .io_maskOut_8_5_1(dataModule_io_maskOut_8_5_1),
    .io_maskOut_8_5_2(dataModule_io_maskOut_8_5_2),
    .io_maskOut_8_5_3(dataModule_io_maskOut_8_5_3),
    .io_maskOut_8_5_4(dataModule_io_maskOut_8_5_4),
    .io_maskOut_8_5_5(dataModule_io_maskOut_8_5_5),
    .io_maskOut_8_5_6(dataModule_io_maskOut_8_5_6),
    .io_maskOut_8_5_7(dataModule_io_maskOut_8_5_7),
    .io_maskOut_8_6_0(dataModule_io_maskOut_8_6_0),
    .io_maskOut_8_6_1(dataModule_io_maskOut_8_6_1),
    .io_maskOut_8_6_2(dataModule_io_maskOut_8_6_2),
    .io_maskOut_8_6_3(dataModule_io_maskOut_8_6_3),
    .io_maskOut_8_6_4(dataModule_io_maskOut_8_6_4),
    .io_maskOut_8_6_5(dataModule_io_maskOut_8_6_5),
    .io_maskOut_8_6_6(dataModule_io_maskOut_8_6_6),
    .io_maskOut_8_6_7(dataModule_io_maskOut_8_6_7),
    .io_maskOut_8_7_0(dataModule_io_maskOut_8_7_0),
    .io_maskOut_8_7_1(dataModule_io_maskOut_8_7_1),
    .io_maskOut_8_7_2(dataModule_io_maskOut_8_7_2),
    .io_maskOut_8_7_3(dataModule_io_maskOut_8_7_3),
    .io_maskOut_8_7_4(dataModule_io_maskOut_8_7_4),
    .io_maskOut_8_7_5(dataModule_io_maskOut_8_7_5),
    .io_maskOut_8_7_6(dataModule_io_maskOut_8_7_6),
    .io_maskOut_8_7_7(dataModule_io_maskOut_8_7_7),
    .io_maskOut_9_0_0(dataModule_io_maskOut_9_0_0),
    .io_maskOut_9_0_1(dataModule_io_maskOut_9_0_1),
    .io_maskOut_9_0_2(dataModule_io_maskOut_9_0_2),
    .io_maskOut_9_0_3(dataModule_io_maskOut_9_0_3),
    .io_maskOut_9_0_4(dataModule_io_maskOut_9_0_4),
    .io_maskOut_9_0_5(dataModule_io_maskOut_9_0_5),
    .io_maskOut_9_0_6(dataModule_io_maskOut_9_0_6),
    .io_maskOut_9_0_7(dataModule_io_maskOut_9_0_7),
    .io_maskOut_9_1_0(dataModule_io_maskOut_9_1_0),
    .io_maskOut_9_1_1(dataModule_io_maskOut_9_1_1),
    .io_maskOut_9_1_2(dataModule_io_maskOut_9_1_2),
    .io_maskOut_9_1_3(dataModule_io_maskOut_9_1_3),
    .io_maskOut_9_1_4(dataModule_io_maskOut_9_1_4),
    .io_maskOut_9_1_5(dataModule_io_maskOut_9_1_5),
    .io_maskOut_9_1_6(dataModule_io_maskOut_9_1_6),
    .io_maskOut_9_1_7(dataModule_io_maskOut_9_1_7),
    .io_maskOut_9_2_0(dataModule_io_maskOut_9_2_0),
    .io_maskOut_9_2_1(dataModule_io_maskOut_9_2_1),
    .io_maskOut_9_2_2(dataModule_io_maskOut_9_2_2),
    .io_maskOut_9_2_3(dataModule_io_maskOut_9_2_3),
    .io_maskOut_9_2_4(dataModule_io_maskOut_9_2_4),
    .io_maskOut_9_2_5(dataModule_io_maskOut_9_2_5),
    .io_maskOut_9_2_6(dataModule_io_maskOut_9_2_6),
    .io_maskOut_9_2_7(dataModule_io_maskOut_9_2_7),
    .io_maskOut_9_3_0(dataModule_io_maskOut_9_3_0),
    .io_maskOut_9_3_1(dataModule_io_maskOut_9_3_1),
    .io_maskOut_9_3_2(dataModule_io_maskOut_9_3_2),
    .io_maskOut_9_3_3(dataModule_io_maskOut_9_3_3),
    .io_maskOut_9_3_4(dataModule_io_maskOut_9_3_4),
    .io_maskOut_9_3_5(dataModule_io_maskOut_9_3_5),
    .io_maskOut_9_3_6(dataModule_io_maskOut_9_3_6),
    .io_maskOut_9_3_7(dataModule_io_maskOut_9_3_7),
    .io_maskOut_9_4_0(dataModule_io_maskOut_9_4_0),
    .io_maskOut_9_4_1(dataModule_io_maskOut_9_4_1),
    .io_maskOut_9_4_2(dataModule_io_maskOut_9_4_2),
    .io_maskOut_9_4_3(dataModule_io_maskOut_9_4_3),
    .io_maskOut_9_4_4(dataModule_io_maskOut_9_4_4),
    .io_maskOut_9_4_5(dataModule_io_maskOut_9_4_5),
    .io_maskOut_9_4_6(dataModule_io_maskOut_9_4_6),
    .io_maskOut_9_4_7(dataModule_io_maskOut_9_4_7),
    .io_maskOut_9_5_0(dataModule_io_maskOut_9_5_0),
    .io_maskOut_9_5_1(dataModule_io_maskOut_9_5_1),
    .io_maskOut_9_5_2(dataModule_io_maskOut_9_5_2),
    .io_maskOut_9_5_3(dataModule_io_maskOut_9_5_3),
    .io_maskOut_9_5_4(dataModule_io_maskOut_9_5_4),
    .io_maskOut_9_5_5(dataModule_io_maskOut_9_5_5),
    .io_maskOut_9_5_6(dataModule_io_maskOut_9_5_6),
    .io_maskOut_9_5_7(dataModule_io_maskOut_9_5_7),
    .io_maskOut_9_6_0(dataModule_io_maskOut_9_6_0),
    .io_maskOut_9_6_1(dataModule_io_maskOut_9_6_1),
    .io_maskOut_9_6_2(dataModule_io_maskOut_9_6_2),
    .io_maskOut_9_6_3(dataModule_io_maskOut_9_6_3),
    .io_maskOut_9_6_4(dataModule_io_maskOut_9_6_4),
    .io_maskOut_9_6_5(dataModule_io_maskOut_9_6_5),
    .io_maskOut_9_6_6(dataModule_io_maskOut_9_6_6),
    .io_maskOut_9_6_7(dataModule_io_maskOut_9_6_7),
    .io_maskOut_9_7_0(dataModule_io_maskOut_9_7_0),
    .io_maskOut_9_7_1(dataModule_io_maskOut_9_7_1),
    .io_maskOut_9_7_2(dataModule_io_maskOut_9_7_2),
    .io_maskOut_9_7_3(dataModule_io_maskOut_9_7_3),
    .io_maskOut_9_7_4(dataModule_io_maskOut_9_7_4),
    .io_maskOut_9_7_5(dataModule_io_maskOut_9_7_5),
    .io_maskOut_9_7_6(dataModule_io_maskOut_9_7_6),
    .io_maskOut_9_7_7(dataModule_io_maskOut_9_7_7),
    .io_maskOut_10_0_0(dataModule_io_maskOut_10_0_0),
    .io_maskOut_10_0_1(dataModule_io_maskOut_10_0_1),
    .io_maskOut_10_0_2(dataModule_io_maskOut_10_0_2),
    .io_maskOut_10_0_3(dataModule_io_maskOut_10_0_3),
    .io_maskOut_10_0_4(dataModule_io_maskOut_10_0_4),
    .io_maskOut_10_0_5(dataModule_io_maskOut_10_0_5),
    .io_maskOut_10_0_6(dataModule_io_maskOut_10_0_6),
    .io_maskOut_10_0_7(dataModule_io_maskOut_10_0_7),
    .io_maskOut_10_1_0(dataModule_io_maskOut_10_1_0),
    .io_maskOut_10_1_1(dataModule_io_maskOut_10_1_1),
    .io_maskOut_10_1_2(dataModule_io_maskOut_10_1_2),
    .io_maskOut_10_1_3(dataModule_io_maskOut_10_1_3),
    .io_maskOut_10_1_4(dataModule_io_maskOut_10_1_4),
    .io_maskOut_10_1_5(dataModule_io_maskOut_10_1_5),
    .io_maskOut_10_1_6(dataModule_io_maskOut_10_1_6),
    .io_maskOut_10_1_7(dataModule_io_maskOut_10_1_7),
    .io_maskOut_10_2_0(dataModule_io_maskOut_10_2_0),
    .io_maskOut_10_2_1(dataModule_io_maskOut_10_2_1),
    .io_maskOut_10_2_2(dataModule_io_maskOut_10_2_2),
    .io_maskOut_10_2_3(dataModule_io_maskOut_10_2_3),
    .io_maskOut_10_2_4(dataModule_io_maskOut_10_2_4),
    .io_maskOut_10_2_5(dataModule_io_maskOut_10_2_5),
    .io_maskOut_10_2_6(dataModule_io_maskOut_10_2_6),
    .io_maskOut_10_2_7(dataModule_io_maskOut_10_2_7),
    .io_maskOut_10_3_0(dataModule_io_maskOut_10_3_0),
    .io_maskOut_10_3_1(dataModule_io_maskOut_10_3_1),
    .io_maskOut_10_3_2(dataModule_io_maskOut_10_3_2),
    .io_maskOut_10_3_3(dataModule_io_maskOut_10_3_3),
    .io_maskOut_10_3_4(dataModule_io_maskOut_10_3_4),
    .io_maskOut_10_3_5(dataModule_io_maskOut_10_3_5),
    .io_maskOut_10_3_6(dataModule_io_maskOut_10_3_6),
    .io_maskOut_10_3_7(dataModule_io_maskOut_10_3_7),
    .io_maskOut_10_4_0(dataModule_io_maskOut_10_4_0),
    .io_maskOut_10_4_1(dataModule_io_maskOut_10_4_1),
    .io_maskOut_10_4_2(dataModule_io_maskOut_10_4_2),
    .io_maskOut_10_4_3(dataModule_io_maskOut_10_4_3),
    .io_maskOut_10_4_4(dataModule_io_maskOut_10_4_4),
    .io_maskOut_10_4_5(dataModule_io_maskOut_10_4_5),
    .io_maskOut_10_4_6(dataModule_io_maskOut_10_4_6),
    .io_maskOut_10_4_7(dataModule_io_maskOut_10_4_7),
    .io_maskOut_10_5_0(dataModule_io_maskOut_10_5_0),
    .io_maskOut_10_5_1(dataModule_io_maskOut_10_5_1),
    .io_maskOut_10_5_2(dataModule_io_maskOut_10_5_2),
    .io_maskOut_10_5_3(dataModule_io_maskOut_10_5_3),
    .io_maskOut_10_5_4(dataModule_io_maskOut_10_5_4),
    .io_maskOut_10_5_5(dataModule_io_maskOut_10_5_5),
    .io_maskOut_10_5_6(dataModule_io_maskOut_10_5_6),
    .io_maskOut_10_5_7(dataModule_io_maskOut_10_5_7),
    .io_maskOut_10_6_0(dataModule_io_maskOut_10_6_0),
    .io_maskOut_10_6_1(dataModule_io_maskOut_10_6_1),
    .io_maskOut_10_6_2(dataModule_io_maskOut_10_6_2),
    .io_maskOut_10_6_3(dataModule_io_maskOut_10_6_3),
    .io_maskOut_10_6_4(dataModule_io_maskOut_10_6_4),
    .io_maskOut_10_6_5(dataModule_io_maskOut_10_6_5),
    .io_maskOut_10_6_6(dataModule_io_maskOut_10_6_6),
    .io_maskOut_10_6_7(dataModule_io_maskOut_10_6_7),
    .io_maskOut_10_7_0(dataModule_io_maskOut_10_7_0),
    .io_maskOut_10_7_1(dataModule_io_maskOut_10_7_1),
    .io_maskOut_10_7_2(dataModule_io_maskOut_10_7_2),
    .io_maskOut_10_7_3(dataModule_io_maskOut_10_7_3),
    .io_maskOut_10_7_4(dataModule_io_maskOut_10_7_4),
    .io_maskOut_10_7_5(dataModule_io_maskOut_10_7_5),
    .io_maskOut_10_7_6(dataModule_io_maskOut_10_7_6),
    .io_maskOut_10_7_7(dataModule_io_maskOut_10_7_7),
    .io_maskOut_11_0_0(dataModule_io_maskOut_11_0_0),
    .io_maskOut_11_0_1(dataModule_io_maskOut_11_0_1),
    .io_maskOut_11_0_2(dataModule_io_maskOut_11_0_2),
    .io_maskOut_11_0_3(dataModule_io_maskOut_11_0_3),
    .io_maskOut_11_0_4(dataModule_io_maskOut_11_0_4),
    .io_maskOut_11_0_5(dataModule_io_maskOut_11_0_5),
    .io_maskOut_11_0_6(dataModule_io_maskOut_11_0_6),
    .io_maskOut_11_0_7(dataModule_io_maskOut_11_0_7),
    .io_maskOut_11_1_0(dataModule_io_maskOut_11_1_0),
    .io_maskOut_11_1_1(dataModule_io_maskOut_11_1_1),
    .io_maskOut_11_1_2(dataModule_io_maskOut_11_1_2),
    .io_maskOut_11_1_3(dataModule_io_maskOut_11_1_3),
    .io_maskOut_11_1_4(dataModule_io_maskOut_11_1_4),
    .io_maskOut_11_1_5(dataModule_io_maskOut_11_1_5),
    .io_maskOut_11_1_6(dataModule_io_maskOut_11_1_6),
    .io_maskOut_11_1_7(dataModule_io_maskOut_11_1_7),
    .io_maskOut_11_2_0(dataModule_io_maskOut_11_2_0),
    .io_maskOut_11_2_1(dataModule_io_maskOut_11_2_1),
    .io_maskOut_11_2_2(dataModule_io_maskOut_11_2_2),
    .io_maskOut_11_2_3(dataModule_io_maskOut_11_2_3),
    .io_maskOut_11_2_4(dataModule_io_maskOut_11_2_4),
    .io_maskOut_11_2_5(dataModule_io_maskOut_11_2_5),
    .io_maskOut_11_2_6(dataModule_io_maskOut_11_2_6),
    .io_maskOut_11_2_7(dataModule_io_maskOut_11_2_7),
    .io_maskOut_11_3_0(dataModule_io_maskOut_11_3_0),
    .io_maskOut_11_3_1(dataModule_io_maskOut_11_3_1),
    .io_maskOut_11_3_2(dataModule_io_maskOut_11_3_2),
    .io_maskOut_11_3_3(dataModule_io_maskOut_11_3_3),
    .io_maskOut_11_3_4(dataModule_io_maskOut_11_3_4),
    .io_maskOut_11_3_5(dataModule_io_maskOut_11_3_5),
    .io_maskOut_11_3_6(dataModule_io_maskOut_11_3_6),
    .io_maskOut_11_3_7(dataModule_io_maskOut_11_3_7),
    .io_maskOut_11_4_0(dataModule_io_maskOut_11_4_0),
    .io_maskOut_11_4_1(dataModule_io_maskOut_11_4_1),
    .io_maskOut_11_4_2(dataModule_io_maskOut_11_4_2),
    .io_maskOut_11_4_3(dataModule_io_maskOut_11_4_3),
    .io_maskOut_11_4_4(dataModule_io_maskOut_11_4_4),
    .io_maskOut_11_4_5(dataModule_io_maskOut_11_4_5),
    .io_maskOut_11_4_6(dataModule_io_maskOut_11_4_6),
    .io_maskOut_11_4_7(dataModule_io_maskOut_11_4_7),
    .io_maskOut_11_5_0(dataModule_io_maskOut_11_5_0),
    .io_maskOut_11_5_1(dataModule_io_maskOut_11_5_1),
    .io_maskOut_11_5_2(dataModule_io_maskOut_11_5_2),
    .io_maskOut_11_5_3(dataModule_io_maskOut_11_5_3),
    .io_maskOut_11_5_4(dataModule_io_maskOut_11_5_4),
    .io_maskOut_11_5_5(dataModule_io_maskOut_11_5_5),
    .io_maskOut_11_5_6(dataModule_io_maskOut_11_5_6),
    .io_maskOut_11_5_7(dataModule_io_maskOut_11_5_7),
    .io_maskOut_11_6_0(dataModule_io_maskOut_11_6_0),
    .io_maskOut_11_6_1(dataModule_io_maskOut_11_6_1),
    .io_maskOut_11_6_2(dataModule_io_maskOut_11_6_2),
    .io_maskOut_11_6_3(dataModule_io_maskOut_11_6_3),
    .io_maskOut_11_6_4(dataModule_io_maskOut_11_6_4),
    .io_maskOut_11_6_5(dataModule_io_maskOut_11_6_5),
    .io_maskOut_11_6_6(dataModule_io_maskOut_11_6_6),
    .io_maskOut_11_6_7(dataModule_io_maskOut_11_6_7),
    .io_maskOut_11_7_0(dataModule_io_maskOut_11_7_0),
    .io_maskOut_11_7_1(dataModule_io_maskOut_11_7_1),
    .io_maskOut_11_7_2(dataModule_io_maskOut_11_7_2),
    .io_maskOut_11_7_3(dataModule_io_maskOut_11_7_3),
    .io_maskOut_11_7_4(dataModule_io_maskOut_11_7_4),
    .io_maskOut_11_7_5(dataModule_io_maskOut_11_7_5),
    .io_maskOut_11_7_6(dataModule_io_maskOut_11_7_6),
    .io_maskOut_11_7_7(dataModule_io_maskOut_11_7_7),
    .io_maskOut_12_0_0(dataModule_io_maskOut_12_0_0),
    .io_maskOut_12_0_1(dataModule_io_maskOut_12_0_1),
    .io_maskOut_12_0_2(dataModule_io_maskOut_12_0_2),
    .io_maskOut_12_0_3(dataModule_io_maskOut_12_0_3),
    .io_maskOut_12_0_4(dataModule_io_maskOut_12_0_4),
    .io_maskOut_12_0_5(dataModule_io_maskOut_12_0_5),
    .io_maskOut_12_0_6(dataModule_io_maskOut_12_0_6),
    .io_maskOut_12_0_7(dataModule_io_maskOut_12_0_7),
    .io_maskOut_12_1_0(dataModule_io_maskOut_12_1_0),
    .io_maskOut_12_1_1(dataModule_io_maskOut_12_1_1),
    .io_maskOut_12_1_2(dataModule_io_maskOut_12_1_2),
    .io_maskOut_12_1_3(dataModule_io_maskOut_12_1_3),
    .io_maskOut_12_1_4(dataModule_io_maskOut_12_1_4),
    .io_maskOut_12_1_5(dataModule_io_maskOut_12_1_5),
    .io_maskOut_12_1_6(dataModule_io_maskOut_12_1_6),
    .io_maskOut_12_1_7(dataModule_io_maskOut_12_1_7),
    .io_maskOut_12_2_0(dataModule_io_maskOut_12_2_0),
    .io_maskOut_12_2_1(dataModule_io_maskOut_12_2_1),
    .io_maskOut_12_2_2(dataModule_io_maskOut_12_2_2),
    .io_maskOut_12_2_3(dataModule_io_maskOut_12_2_3),
    .io_maskOut_12_2_4(dataModule_io_maskOut_12_2_4),
    .io_maskOut_12_2_5(dataModule_io_maskOut_12_2_5),
    .io_maskOut_12_2_6(dataModule_io_maskOut_12_2_6),
    .io_maskOut_12_2_7(dataModule_io_maskOut_12_2_7),
    .io_maskOut_12_3_0(dataModule_io_maskOut_12_3_0),
    .io_maskOut_12_3_1(dataModule_io_maskOut_12_3_1),
    .io_maskOut_12_3_2(dataModule_io_maskOut_12_3_2),
    .io_maskOut_12_3_3(dataModule_io_maskOut_12_3_3),
    .io_maskOut_12_3_4(dataModule_io_maskOut_12_3_4),
    .io_maskOut_12_3_5(dataModule_io_maskOut_12_3_5),
    .io_maskOut_12_3_6(dataModule_io_maskOut_12_3_6),
    .io_maskOut_12_3_7(dataModule_io_maskOut_12_3_7),
    .io_maskOut_12_4_0(dataModule_io_maskOut_12_4_0),
    .io_maskOut_12_4_1(dataModule_io_maskOut_12_4_1),
    .io_maskOut_12_4_2(dataModule_io_maskOut_12_4_2),
    .io_maskOut_12_4_3(dataModule_io_maskOut_12_4_3),
    .io_maskOut_12_4_4(dataModule_io_maskOut_12_4_4),
    .io_maskOut_12_4_5(dataModule_io_maskOut_12_4_5),
    .io_maskOut_12_4_6(dataModule_io_maskOut_12_4_6),
    .io_maskOut_12_4_7(dataModule_io_maskOut_12_4_7),
    .io_maskOut_12_5_0(dataModule_io_maskOut_12_5_0),
    .io_maskOut_12_5_1(dataModule_io_maskOut_12_5_1),
    .io_maskOut_12_5_2(dataModule_io_maskOut_12_5_2),
    .io_maskOut_12_5_3(dataModule_io_maskOut_12_5_3),
    .io_maskOut_12_5_4(dataModule_io_maskOut_12_5_4),
    .io_maskOut_12_5_5(dataModule_io_maskOut_12_5_5),
    .io_maskOut_12_5_6(dataModule_io_maskOut_12_5_6),
    .io_maskOut_12_5_7(dataModule_io_maskOut_12_5_7),
    .io_maskOut_12_6_0(dataModule_io_maskOut_12_6_0),
    .io_maskOut_12_6_1(dataModule_io_maskOut_12_6_1),
    .io_maskOut_12_6_2(dataModule_io_maskOut_12_6_2),
    .io_maskOut_12_6_3(dataModule_io_maskOut_12_6_3),
    .io_maskOut_12_6_4(dataModule_io_maskOut_12_6_4),
    .io_maskOut_12_6_5(dataModule_io_maskOut_12_6_5),
    .io_maskOut_12_6_6(dataModule_io_maskOut_12_6_6),
    .io_maskOut_12_6_7(dataModule_io_maskOut_12_6_7),
    .io_maskOut_12_7_0(dataModule_io_maskOut_12_7_0),
    .io_maskOut_12_7_1(dataModule_io_maskOut_12_7_1),
    .io_maskOut_12_7_2(dataModule_io_maskOut_12_7_2),
    .io_maskOut_12_7_3(dataModule_io_maskOut_12_7_3),
    .io_maskOut_12_7_4(dataModule_io_maskOut_12_7_4),
    .io_maskOut_12_7_5(dataModule_io_maskOut_12_7_5),
    .io_maskOut_12_7_6(dataModule_io_maskOut_12_7_6),
    .io_maskOut_12_7_7(dataModule_io_maskOut_12_7_7),
    .io_maskOut_13_0_0(dataModule_io_maskOut_13_0_0),
    .io_maskOut_13_0_1(dataModule_io_maskOut_13_0_1),
    .io_maskOut_13_0_2(dataModule_io_maskOut_13_0_2),
    .io_maskOut_13_0_3(dataModule_io_maskOut_13_0_3),
    .io_maskOut_13_0_4(dataModule_io_maskOut_13_0_4),
    .io_maskOut_13_0_5(dataModule_io_maskOut_13_0_5),
    .io_maskOut_13_0_6(dataModule_io_maskOut_13_0_6),
    .io_maskOut_13_0_7(dataModule_io_maskOut_13_0_7),
    .io_maskOut_13_1_0(dataModule_io_maskOut_13_1_0),
    .io_maskOut_13_1_1(dataModule_io_maskOut_13_1_1),
    .io_maskOut_13_1_2(dataModule_io_maskOut_13_1_2),
    .io_maskOut_13_1_3(dataModule_io_maskOut_13_1_3),
    .io_maskOut_13_1_4(dataModule_io_maskOut_13_1_4),
    .io_maskOut_13_1_5(dataModule_io_maskOut_13_1_5),
    .io_maskOut_13_1_6(dataModule_io_maskOut_13_1_6),
    .io_maskOut_13_1_7(dataModule_io_maskOut_13_1_7),
    .io_maskOut_13_2_0(dataModule_io_maskOut_13_2_0),
    .io_maskOut_13_2_1(dataModule_io_maskOut_13_2_1),
    .io_maskOut_13_2_2(dataModule_io_maskOut_13_2_2),
    .io_maskOut_13_2_3(dataModule_io_maskOut_13_2_3),
    .io_maskOut_13_2_4(dataModule_io_maskOut_13_2_4),
    .io_maskOut_13_2_5(dataModule_io_maskOut_13_2_5),
    .io_maskOut_13_2_6(dataModule_io_maskOut_13_2_6),
    .io_maskOut_13_2_7(dataModule_io_maskOut_13_2_7),
    .io_maskOut_13_3_0(dataModule_io_maskOut_13_3_0),
    .io_maskOut_13_3_1(dataModule_io_maskOut_13_3_1),
    .io_maskOut_13_3_2(dataModule_io_maskOut_13_3_2),
    .io_maskOut_13_3_3(dataModule_io_maskOut_13_3_3),
    .io_maskOut_13_3_4(dataModule_io_maskOut_13_3_4),
    .io_maskOut_13_3_5(dataModule_io_maskOut_13_3_5),
    .io_maskOut_13_3_6(dataModule_io_maskOut_13_3_6),
    .io_maskOut_13_3_7(dataModule_io_maskOut_13_3_7),
    .io_maskOut_13_4_0(dataModule_io_maskOut_13_4_0),
    .io_maskOut_13_4_1(dataModule_io_maskOut_13_4_1),
    .io_maskOut_13_4_2(dataModule_io_maskOut_13_4_2),
    .io_maskOut_13_4_3(dataModule_io_maskOut_13_4_3),
    .io_maskOut_13_4_4(dataModule_io_maskOut_13_4_4),
    .io_maskOut_13_4_5(dataModule_io_maskOut_13_4_5),
    .io_maskOut_13_4_6(dataModule_io_maskOut_13_4_6),
    .io_maskOut_13_4_7(dataModule_io_maskOut_13_4_7),
    .io_maskOut_13_5_0(dataModule_io_maskOut_13_5_0),
    .io_maskOut_13_5_1(dataModule_io_maskOut_13_5_1),
    .io_maskOut_13_5_2(dataModule_io_maskOut_13_5_2),
    .io_maskOut_13_5_3(dataModule_io_maskOut_13_5_3),
    .io_maskOut_13_5_4(dataModule_io_maskOut_13_5_4),
    .io_maskOut_13_5_5(dataModule_io_maskOut_13_5_5),
    .io_maskOut_13_5_6(dataModule_io_maskOut_13_5_6),
    .io_maskOut_13_5_7(dataModule_io_maskOut_13_5_7),
    .io_maskOut_13_6_0(dataModule_io_maskOut_13_6_0),
    .io_maskOut_13_6_1(dataModule_io_maskOut_13_6_1),
    .io_maskOut_13_6_2(dataModule_io_maskOut_13_6_2),
    .io_maskOut_13_6_3(dataModule_io_maskOut_13_6_3),
    .io_maskOut_13_6_4(dataModule_io_maskOut_13_6_4),
    .io_maskOut_13_6_5(dataModule_io_maskOut_13_6_5),
    .io_maskOut_13_6_6(dataModule_io_maskOut_13_6_6),
    .io_maskOut_13_6_7(dataModule_io_maskOut_13_6_7),
    .io_maskOut_13_7_0(dataModule_io_maskOut_13_7_0),
    .io_maskOut_13_7_1(dataModule_io_maskOut_13_7_1),
    .io_maskOut_13_7_2(dataModule_io_maskOut_13_7_2),
    .io_maskOut_13_7_3(dataModule_io_maskOut_13_7_3),
    .io_maskOut_13_7_4(dataModule_io_maskOut_13_7_4),
    .io_maskOut_13_7_5(dataModule_io_maskOut_13_7_5),
    .io_maskOut_13_7_6(dataModule_io_maskOut_13_7_6),
    .io_maskOut_13_7_7(dataModule_io_maskOut_13_7_7),
    .io_maskOut_14_0_0(dataModule_io_maskOut_14_0_0),
    .io_maskOut_14_0_1(dataModule_io_maskOut_14_0_1),
    .io_maskOut_14_0_2(dataModule_io_maskOut_14_0_2),
    .io_maskOut_14_0_3(dataModule_io_maskOut_14_0_3),
    .io_maskOut_14_0_4(dataModule_io_maskOut_14_0_4),
    .io_maskOut_14_0_5(dataModule_io_maskOut_14_0_5),
    .io_maskOut_14_0_6(dataModule_io_maskOut_14_0_6),
    .io_maskOut_14_0_7(dataModule_io_maskOut_14_0_7),
    .io_maskOut_14_1_0(dataModule_io_maskOut_14_1_0),
    .io_maskOut_14_1_1(dataModule_io_maskOut_14_1_1),
    .io_maskOut_14_1_2(dataModule_io_maskOut_14_1_2),
    .io_maskOut_14_1_3(dataModule_io_maskOut_14_1_3),
    .io_maskOut_14_1_4(dataModule_io_maskOut_14_1_4),
    .io_maskOut_14_1_5(dataModule_io_maskOut_14_1_5),
    .io_maskOut_14_1_6(dataModule_io_maskOut_14_1_6),
    .io_maskOut_14_1_7(dataModule_io_maskOut_14_1_7),
    .io_maskOut_14_2_0(dataModule_io_maskOut_14_2_0),
    .io_maskOut_14_2_1(dataModule_io_maskOut_14_2_1),
    .io_maskOut_14_2_2(dataModule_io_maskOut_14_2_2),
    .io_maskOut_14_2_3(dataModule_io_maskOut_14_2_3),
    .io_maskOut_14_2_4(dataModule_io_maskOut_14_2_4),
    .io_maskOut_14_2_5(dataModule_io_maskOut_14_2_5),
    .io_maskOut_14_2_6(dataModule_io_maskOut_14_2_6),
    .io_maskOut_14_2_7(dataModule_io_maskOut_14_2_7),
    .io_maskOut_14_3_0(dataModule_io_maskOut_14_3_0),
    .io_maskOut_14_3_1(dataModule_io_maskOut_14_3_1),
    .io_maskOut_14_3_2(dataModule_io_maskOut_14_3_2),
    .io_maskOut_14_3_3(dataModule_io_maskOut_14_3_3),
    .io_maskOut_14_3_4(dataModule_io_maskOut_14_3_4),
    .io_maskOut_14_3_5(dataModule_io_maskOut_14_3_5),
    .io_maskOut_14_3_6(dataModule_io_maskOut_14_3_6),
    .io_maskOut_14_3_7(dataModule_io_maskOut_14_3_7),
    .io_maskOut_14_4_0(dataModule_io_maskOut_14_4_0),
    .io_maskOut_14_4_1(dataModule_io_maskOut_14_4_1),
    .io_maskOut_14_4_2(dataModule_io_maskOut_14_4_2),
    .io_maskOut_14_4_3(dataModule_io_maskOut_14_4_3),
    .io_maskOut_14_4_4(dataModule_io_maskOut_14_4_4),
    .io_maskOut_14_4_5(dataModule_io_maskOut_14_4_5),
    .io_maskOut_14_4_6(dataModule_io_maskOut_14_4_6),
    .io_maskOut_14_4_7(dataModule_io_maskOut_14_4_7),
    .io_maskOut_14_5_0(dataModule_io_maskOut_14_5_0),
    .io_maskOut_14_5_1(dataModule_io_maskOut_14_5_1),
    .io_maskOut_14_5_2(dataModule_io_maskOut_14_5_2),
    .io_maskOut_14_5_3(dataModule_io_maskOut_14_5_3),
    .io_maskOut_14_5_4(dataModule_io_maskOut_14_5_4),
    .io_maskOut_14_5_5(dataModule_io_maskOut_14_5_5),
    .io_maskOut_14_5_6(dataModule_io_maskOut_14_5_6),
    .io_maskOut_14_5_7(dataModule_io_maskOut_14_5_7),
    .io_maskOut_14_6_0(dataModule_io_maskOut_14_6_0),
    .io_maskOut_14_6_1(dataModule_io_maskOut_14_6_1),
    .io_maskOut_14_6_2(dataModule_io_maskOut_14_6_2),
    .io_maskOut_14_6_3(dataModule_io_maskOut_14_6_3),
    .io_maskOut_14_6_4(dataModule_io_maskOut_14_6_4),
    .io_maskOut_14_6_5(dataModule_io_maskOut_14_6_5),
    .io_maskOut_14_6_6(dataModule_io_maskOut_14_6_6),
    .io_maskOut_14_6_7(dataModule_io_maskOut_14_6_7),
    .io_maskOut_14_7_0(dataModule_io_maskOut_14_7_0),
    .io_maskOut_14_7_1(dataModule_io_maskOut_14_7_1),
    .io_maskOut_14_7_2(dataModule_io_maskOut_14_7_2),
    .io_maskOut_14_7_3(dataModule_io_maskOut_14_7_3),
    .io_maskOut_14_7_4(dataModule_io_maskOut_14_7_4),
    .io_maskOut_14_7_5(dataModule_io_maskOut_14_7_5),
    .io_maskOut_14_7_6(dataModule_io_maskOut_14_7_6),
    .io_maskOut_14_7_7(dataModule_io_maskOut_14_7_7),
    .io_maskOut_15_0_0(dataModule_io_maskOut_15_0_0),
    .io_maskOut_15_0_1(dataModule_io_maskOut_15_0_1),
    .io_maskOut_15_0_2(dataModule_io_maskOut_15_0_2),
    .io_maskOut_15_0_3(dataModule_io_maskOut_15_0_3),
    .io_maskOut_15_0_4(dataModule_io_maskOut_15_0_4),
    .io_maskOut_15_0_5(dataModule_io_maskOut_15_0_5),
    .io_maskOut_15_0_6(dataModule_io_maskOut_15_0_6),
    .io_maskOut_15_0_7(dataModule_io_maskOut_15_0_7),
    .io_maskOut_15_1_0(dataModule_io_maskOut_15_1_0),
    .io_maskOut_15_1_1(dataModule_io_maskOut_15_1_1),
    .io_maskOut_15_1_2(dataModule_io_maskOut_15_1_2),
    .io_maskOut_15_1_3(dataModule_io_maskOut_15_1_3),
    .io_maskOut_15_1_4(dataModule_io_maskOut_15_1_4),
    .io_maskOut_15_1_5(dataModule_io_maskOut_15_1_5),
    .io_maskOut_15_1_6(dataModule_io_maskOut_15_1_6),
    .io_maskOut_15_1_7(dataModule_io_maskOut_15_1_7),
    .io_maskOut_15_2_0(dataModule_io_maskOut_15_2_0),
    .io_maskOut_15_2_1(dataModule_io_maskOut_15_2_1),
    .io_maskOut_15_2_2(dataModule_io_maskOut_15_2_2),
    .io_maskOut_15_2_3(dataModule_io_maskOut_15_2_3),
    .io_maskOut_15_2_4(dataModule_io_maskOut_15_2_4),
    .io_maskOut_15_2_5(dataModule_io_maskOut_15_2_5),
    .io_maskOut_15_2_6(dataModule_io_maskOut_15_2_6),
    .io_maskOut_15_2_7(dataModule_io_maskOut_15_2_7),
    .io_maskOut_15_3_0(dataModule_io_maskOut_15_3_0),
    .io_maskOut_15_3_1(dataModule_io_maskOut_15_3_1),
    .io_maskOut_15_3_2(dataModule_io_maskOut_15_3_2),
    .io_maskOut_15_3_3(dataModule_io_maskOut_15_3_3),
    .io_maskOut_15_3_4(dataModule_io_maskOut_15_3_4),
    .io_maskOut_15_3_5(dataModule_io_maskOut_15_3_5),
    .io_maskOut_15_3_6(dataModule_io_maskOut_15_3_6),
    .io_maskOut_15_3_7(dataModule_io_maskOut_15_3_7),
    .io_maskOut_15_4_0(dataModule_io_maskOut_15_4_0),
    .io_maskOut_15_4_1(dataModule_io_maskOut_15_4_1),
    .io_maskOut_15_4_2(dataModule_io_maskOut_15_4_2),
    .io_maskOut_15_4_3(dataModule_io_maskOut_15_4_3),
    .io_maskOut_15_4_4(dataModule_io_maskOut_15_4_4),
    .io_maskOut_15_4_5(dataModule_io_maskOut_15_4_5),
    .io_maskOut_15_4_6(dataModule_io_maskOut_15_4_6),
    .io_maskOut_15_4_7(dataModule_io_maskOut_15_4_7),
    .io_maskOut_15_5_0(dataModule_io_maskOut_15_5_0),
    .io_maskOut_15_5_1(dataModule_io_maskOut_15_5_1),
    .io_maskOut_15_5_2(dataModule_io_maskOut_15_5_2),
    .io_maskOut_15_5_3(dataModule_io_maskOut_15_5_3),
    .io_maskOut_15_5_4(dataModule_io_maskOut_15_5_4),
    .io_maskOut_15_5_5(dataModule_io_maskOut_15_5_5),
    .io_maskOut_15_5_6(dataModule_io_maskOut_15_5_6),
    .io_maskOut_15_5_7(dataModule_io_maskOut_15_5_7),
    .io_maskOut_15_6_0(dataModule_io_maskOut_15_6_0),
    .io_maskOut_15_6_1(dataModule_io_maskOut_15_6_1),
    .io_maskOut_15_6_2(dataModule_io_maskOut_15_6_2),
    .io_maskOut_15_6_3(dataModule_io_maskOut_15_6_3),
    .io_maskOut_15_6_4(dataModule_io_maskOut_15_6_4),
    .io_maskOut_15_6_5(dataModule_io_maskOut_15_6_5),
    .io_maskOut_15_6_6(dataModule_io_maskOut_15_6_6),
    .io_maskOut_15_6_7(dataModule_io_maskOut_15_6_7),
    .io_maskOut_15_7_0(dataModule_io_maskOut_15_7_0),
    .io_maskOut_15_7_1(dataModule_io_maskOut_15_7_1),
    .io_maskOut_15_7_2(dataModule_io_maskOut_15_7_2),
    .io_maskOut_15_7_3(dataModule_io_maskOut_15_7_3),
    .io_maskOut_15_7_4(dataModule_io_maskOut_15_7_4),
    .io_maskOut_15_7_5(dataModule_io_maskOut_15_7_5),
    .io_maskOut_15_7_6(dataModule_io_maskOut_15_7_6),
    .io_maskOut_15_7_7(dataModule_io_maskOut_15_7_7)
  );
  ValidPLRUWrapper Sbuffer_PLRU ( // @[Sbuffer.scala 324:20]
    .clock(Sbuffer_PLRU_clock),
    .reset(Sbuffer_PLRU_reset),
    .io_access_0_valid(Sbuffer_PLRU_io_access_0_valid),
    .io_access_0_bits(Sbuffer_PLRU_io_access_0_bits),
    .io_access_1_valid(Sbuffer_PLRU_io_access_1_valid),
    .io_access_1_bits(Sbuffer_PLRU_io_access_1_bits),
    .io_access_2_valid(Sbuffer_PLRU_io_access_2_valid),
    .io_access_2_bits(Sbuffer_PLRU_io_access_2_bits),
    .io_candidateVec_0(Sbuffer_PLRU_io_candidateVec_0),
    .io_candidateVec_1(Sbuffer_PLRU_io_candidateVec_1),
    .io_candidateVec_2(Sbuffer_PLRU_io_candidateVec_2),
    .io_candidateVec_3(Sbuffer_PLRU_io_candidateVec_3),
    .io_candidateVec_4(Sbuffer_PLRU_io_candidateVec_4),
    .io_candidateVec_5(Sbuffer_PLRU_io_candidateVec_5),
    .io_candidateVec_6(Sbuffer_PLRU_io_candidateVec_6),
    .io_candidateVec_7(Sbuffer_PLRU_io_candidateVec_7),
    .io_candidateVec_8(Sbuffer_PLRU_io_candidateVec_8),
    .io_candidateVec_9(Sbuffer_PLRU_io_candidateVec_9),
    .io_candidateVec_10(Sbuffer_PLRU_io_candidateVec_10),
    .io_candidateVec_11(Sbuffer_PLRU_io_candidateVec_11),
    .io_candidateVec_12(Sbuffer_PLRU_io_candidateVec_12),
    .io_candidateVec_13(Sbuffer_PLRU_io_candidateVec_13),
    .io_candidateVec_14(Sbuffer_PLRU_io_candidateVec_14),
    .io_candidateVec_15(Sbuffer_PLRU_io_candidateVec_15),
    .io_replaceWay(Sbuffer_PLRU_io_replaceWay)
  );
  assign io_in_0_ready = sbuffer_state != 2'h3 & _firstCanInsert_T_1; // @[Sbuffer.scala 434:58]
  assign io_in_1_ready = secondCanInsert & ~sameWord & io_in_0_ready; // @[Sbuffer.scala 445:50]
  assign io_dcache_req_valid = sbuffer_out_s1_valid & _sbuffer_out_s1_ready_T; // @[Sbuffer.scala 698:47]
  assign io_dcache_req_bits_vaddr = {sbuffer_out_s1_evictionVTag,6'h0}; // @[Cat.scala 33:92]
  assign io_dcache_req_bits_addr = {sbuffer_out_s1_evictionPTag,6'h0}; // @[Cat.scala 33:92]
  assign io_dcache_req_bits_data = {io_dcache_req_bits_data_hi,io_dcache_req_bits_data_lo}; // @[Sbuffer.scala 703:64]
  assign io_dcache_req_bits_mask = {io_dcache_req_bits_mask_hi,io_dcache_req_bits_mask_lo}; // @[Sbuffer.scala 704:64]
  assign io_dcache_req_bits_id = {{2'd0}, sbuffer_out_s1_evictionIdx}; // @[Sbuffer.scala 705:25]
  assign io_forward_0_forwardMask_0 = selectedValidMask_0_0 | selectedInflightMask_0_0; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_1 = selectedValidMask_0_1 | selectedInflightMask_0_1; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_2 = selectedValidMask_0_2 | selectedInflightMask_0_2; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_3 = selectedValidMask_0_3 | selectedInflightMask_0_3; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_4 = selectedValidMask_0_4 | selectedInflightMask_0_4; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_5 = selectedValidMask_0_5 | selectedInflightMask_0_5; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_6 = selectedValidMask_0_6 | selectedInflightMask_0_6; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardMask_7 = selectedValidMask_0_7 | selectedInflightMask_0_7; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_0_forwardData_0 = selectedValidMask_0_0 ? selectedValidData_0_0 : selectedInflightData_0_0; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_1 = selectedValidMask_0_1 ? selectedValidData_0_1 : selectedInflightData_0_1; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_2 = selectedValidMask_0_2 ? selectedValidData_0_2 : selectedInflightData_0_2; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_3 = selectedValidMask_0_3 ? selectedValidData_0_3 : selectedInflightData_0_3; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_4 = selectedValidMask_0_4 ? selectedValidData_0_4 : selectedInflightData_0_4; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_5 = selectedValidMask_0_5 ? selectedValidData_0_5 : selectedInflightData_0_5; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_6 = selectedValidMask_0_6 ? selectedValidData_0_6 : selectedInflightData_0_6; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_forwardData_7 = selectedValidMask_0_7 ? selectedValidData_0_7 : selectedInflightData_0_7; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_0_matchInvalid = tag_mismatch_REG & _tag_mismatch_T_49; // @[Sbuffer.scala 799:47]
  assign io_forward_1_forwardMask_0 = selectedValidMask_1_0 | selectedInflightMask_1_0; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_1 = selectedValidMask_1_1 | selectedInflightMask_1_1; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_2 = selectedValidMask_1_2 | selectedInflightMask_1_2; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_3 = selectedValidMask_1_3 | selectedInflightMask_1_3; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_4 = selectedValidMask_1_4 | selectedInflightMask_1_4; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_5 = selectedValidMask_1_5 | selectedInflightMask_1_5; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_6 = selectedValidMask_1_6 | selectedInflightMask_1_6; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardMask_7 = selectedValidMask_1_7 | selectedInflightMask_1_7; // @[Sbuffer.scala 853:34 854:32]
  assign io_forward_1_forwardData_0 = selectedValidMask_1_0 ? selectedValidData_1_0 : selectedInflightData_1_0; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_1 = selectedValidMask_1_1 ? selectedValidData_1_1 : selectedInflightData_1_1; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_2 = selectedValidMask_1_2 ? selectedValidData_1_2 : selectedInflightData_1_2; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_3 = selectedValidMask_1_3 ? selectedValidData_1_3 : selectedInflightData_1_3; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_4 = selectedValidMask_1_4 ? selectedValidData_1_4 : selectedInflightData_1_4; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_5 = selectedValidMask_1_5 ? selectedValidData_1_5 : selectedInflightData_1_5; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_6 = selectedValidMask_1_6 ? selectedValidData_1_6 : selectedInflightData_1_6; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_forwardData_7 = selectedValidMask_1_7 ? selectedValidData_1_7 : selectedInflightData_1_7; // @[Sbuffer.scala 853:34 855:32]
  assign io_forward_1_matchInvalid = tag_mismatch_REG_33 & _tag_mismatch_T_99; // @[Sbuffer.scala 799:47]
  assign io_flush_empty = io_flush_empty_REG; // @[Sbuffer.scala 557:18]
  assign io_perf_0_value = {{4'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_1_value = {{4'd0}, io_perf_1_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_2_value = {{4'd0}, io_perf_2_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_3_value = {{4'd0}, io_perf_3_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_4_value = {{5'd0}, io_perf_4_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_5_value = {{5'd0}, io_perf_5_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_6_value = {{5'd0}, io_perf_6_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_7_value = {{5'd0}, io_perf_7_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_8_value = {{5'd0}, io_perf_8_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_9_value = {{5'd0}, io_perf_9_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_10_value = {{5'd0}, io_perf_10_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_11_value = {{5'd0}, io_perf_11_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_12_value = {{5'd0}, io_perf_12_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_13_value = {{5'd0}, io_perf_13_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_14_value = {{5'd0}, io_perf_14_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_15_value = {{5'd0}, io_perf_15_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign io_perf_16_value = {{5'd0}, io_perf_16_value_REG_1}; // @[PerfCounterUtils.scala 172:17]
  assign dataModule_clock = clock;
  assign dataModule_reset = reset;
  assign dataModule_io_writeReq_0_valid = io_in_0_ready & io_in_0_valid; // @[Decoupled.scala 51:35]
  assign dataModule_io_writeReq_0_bits_wvec = canMerge_0 ? mergeVec_0 : firstInsertVec; // @[Sbuffer.scala 512:24 513:31 517:31]
  assign dataModule_io_writeReq_0_bits_mask = io_in_0_bits_mask; // @[Sbuffer.scala 502:27]
  assign dataModule_io_writeReq_0_bits_data = io_in_0_bits_data; // @[Sbuffer.scala 503:27]
  assign dataModule_io_writeReq_0_bits_wordOffset = io_in_0_bits_addr[35:3]; // @[Sbuffer.scala 306:7]
  assign dataModule_io_writeReq_0_bits_wline = io_in_0_bits_wline; // @[Sbuffer.scala 504:28]
  assign dataModule_io_writeReq_1_valid = io_in_1_ready & io_in_1_valid; // @[Decoupled.scala 51:35]
  assign dataModule_io_writeReq_1_bits_wvec = canMerge_1 ? mergeVec_1 : secondInsertVec; // @[Sbuffer.scala 512:24 513:31 517:31]
  assign dataModule_io_writeReq_1_bits_mask = io_in_1_bits_mask; // @[Sbuffer.scala 502:27]
  assign dataModule_io_writeReq_1_bits_data = io_in_1_bits_data; // @[Sbuffer.scala 503:27]
  assign dataModule_io_writeReq_1_bits_wordOffset = io_in_1_bits_addr[35:3]; // @[Sbuffer.scala 306:7]
  assign dataModule_io_writeReq_1_bits_wline = io_in_1_bits_wline; // @[Sbuffer.scala 504:28]
  assign dataModule_io_maskFlushReq_0_valid = io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 752:21]
  assign dataModule_io_maskFlushReq_0_bits_wvec = _dataModule_io_maskFlushReq_0_bits_wvec_T[15:0]; // @[Sbuffer.scala 753:25]
  assign dataModule_io_maskFlushReq_1_valid = io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 752:21]
  assign dataModule_io_maskFlushReq_1_bits_wvec = _dataModule_io_maskFlushReq_1_bits_wvec_T[15:0]; // @[Sbuffer.scala 753:25]
  assign Sbuffer_PLRU_clock = clock;
  assign Sbuffer_PLRU_reset = reset;
  assign Sbuffer_PLRU_io_access_0_valid = accessIdx_0_valid_REG; // @[Sbuffer.scala 327:23 509:24]
  assign Sbuffer_PLRU_io_access_0_bits = accessIdx_0_bits_REG; // @[Sbuffer.scala 327:23 510:23]
  assign Sbuffer_PLRU_io_access_1_valid = accessIdx_1_valid_REG; // @[Sbuffer.scala 327:23 509:24]
  assign Sbuffer_PLRU_io_access_1_bits = accessIdx_1_bits_REG; // @[Sbuffer.scala 327:23 510:23]
  assign Sbuffer_PLRU_io_access_2_valid = _GEN_888 | _accessIdx_2_valid_T_7; // @[Sbuffer.scala 691:62]
  assign Sbuffer_PLRU_io_access_2_bits = Sbuffer_PLRU_io_replaceWay; // @[Sbuffer.scala 327:23 693:34]
  assign Sbuffer_PLRU_io_candidateVec_0 = stateVec_0_state_valid & ~stateVec_0_state_inflight & ~
    stateVec_0_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_1 = stateVec_1_state_valid & ~stateVec_1_state_inflight & ~
    stateVec_1_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_2 = stateVec_2_state_valid & ~stateVec_2_state_inflight & ~
    stateVec_2_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_3 = stateVec_3_state_valid & ~stateVec_3_state_inflight & ~
    stateVec_3_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_4 = stateVec_4_state_valid & ~stateVec_4_state_inflight & ~
    stateVec_4_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_5 = stateVec_5_state_valid & ~stateVec_5_state_inflight & ~
    stateVec_5_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_6 = stateVec_6_state_valid & ~stateVec_6_state_inflight & ~
    stateVec_6_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_7 = stateVec_7_state_valid & ~stateVec_7_state_inflight & ~
    stateVec_7_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_8 = stateVec_8_state_valid & ~stateVec_8_state_inflight & ~
    stateVec_8_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_9 = stateVec_9_state_valid & ~stateVec_9_state_inflight & ~
    stateVec_9_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_10 = stateVec_10_state_valid & ~stateVec_10_state_inflight & ~
    stateVec_10_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_11 = stateVec_11_state_valid & ~stateVec_11_state_inflight & ~
    stateVec_11_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_12 = stateVec_12_state_valid & ~stateVec_12_state_inflight & ~
    stateVec_12_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_13 = stateVec_13_state_valid & ~stateVec_13_state_inflight & ~
    stateVec_13_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_14 = stateVec_14_state_valid & ~stateVec_14_state_inflight & ~
    stateVec_14_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  assign Sbuffer_PLRU_io_candidateVec_15 = stateVec_15_state_valid & ~stateVec_15_state_inflight & ~
    stateVec_15_w_sameblock_inflight; // @[Sbuffer.scala 66:69]
  always @(posedge clock) begin
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_0 <= _GEN_281;
      end else if (secondInsertVec[0]) begin // @[Sbuffer.scala 458:32]
        ptag_0 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_0 <= _GEN_281;
      end
    end else begin
      ptag_0 <= _GEN_281;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_1 <= _GEN_286;
      end else if (secondInsertVec[1]) begin // @[Sbuffer.scala 458:32]
        ptag_1 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_1 <= _GEN_286;
      end
    end else begin
      ptag_1 <= _GEN_286;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_2 <= _GEN_291;
      end else if (secondInsertVec[2]) begin // @[Sbuffer.scala 458:32]
        ptag_2 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_2 <= _GEN_291;
      end
    end else begin
      ptag_2 <= _GEN_291;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_3 <= _GEN_296;
      end else if (secondInsertVec[3]) begin // @[Sbuffer.scala 458:32]
        ptag_3 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_3 <= _GEN_296;
      end
    end else begin
      ptag_3 <= _GEN_296;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_4 <= _GEN_301;
      end else if (secondInsertVec[4]) begin // @[Sbuffer.scala 458:32]
        ptag_4 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_4 <= _GEN_301;
      end
    end else begin
      ptag_4 <= _GEN_301;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_5 <= _GEN_306;
      end else if (secondInsertVec[5]) begin // @[Sbuffer.scala 458:32]
        ptag_5 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_5 <= _GEN_306;
      end
    end else begin
      ptag_5 <= _GEN_306;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_6 <= _GEN_311;
      end else if (secondInsertVec[6]) begin // @[Sbuffer.scala 458:32]
        ptag_6 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_6 <= _GEN_311;
      end
    end else begin
      ptag_6 <= _GEN_311;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_7 <= _GEN_316;
      end else if (secondInsertVec[7]) begin // @[Sbuffer.scala 458:32]
        ptag_7 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_7 <= _GEN_316;
      end
    end else begin
      ptag_7 <= _GEN_316;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_8 <= _GEN_321;
      end else if (secondInsertVec[8]) begin // @[Sbuffer.scala 458:32]
        ptag_8 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_8 <= _GEN_321;
      end
    end else begin
      ptag_8 <= _GEN_321;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_9 <= _GEN_326;
      end else if (secondInsertVec[9]) begin // @[Sbuffer.scala 458:32]
        ptag_9 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_9 <= _GEN_326;
      end
    end else begin
      ptag_9 <= _GEN_326;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_10 <= _GEN_331;
      end else if (secondInsertVec[10]) begin // @[Sbuffer.scala 458:32]
        ptag_10 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_10 <= _GEN_331;
      end
    end else begin
      ptag_10 <= _GEN_331;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_11 <= _GEN_336;
      end else if (secondInsertVec[11]) begin // @[Sbuffer.scala 458:32]
        ptag_11 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_11 <= _GEN_336;
      end
    end else begin
      ptag_11 <= _GEN_336;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_12 <= _GEN_341;
      end else if (secondInsertVec[12]) begin // @[Sbuffer.scala 458:32]
        ptag_12 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_12 <= _GEN_341;
      end
    end else begin
      ptag_12 <= _GEN_341;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_13 <= _GEN_346;
      end else if (secondInsertVec[13]) begin // @[Sbuffer.scala 458:32]
        ptag_13 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_13 <= _GEN_346;
      end
    end else begin
      ptag_13 <= _GEN_346;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_14 <= _GEN_351;
      end else if (secondInsertVec[14]) begin // @[Sbuffer.scala 458:32]
        ptag_14 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_14 <= _GEN_351;
      end
    end else begin
      ptag_14 <= _GEN_351;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        ptag_15 <= _GEN_356;
      end else if (secondInsertVec[15]) begin // @[Sbuffer.scala 458:32]
        ptag_15 <= inptags_1; // @[Sbuffer.scala 466:24]
      end else begin
        ptag_15 <= _GEN_356;
      end
    end else begin
      ptag_15 <= _GEN_356;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_0 <= _GEN_282;
      end else if (secondInsertVec[0]) begin // @[Sbuffer.scala 458:32]
        vtag_0 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_0 <= _GEN_282;
      end
    end else begin
      vtag_0 <= _GEN_282;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_1 <= _GEN_287;
      end else if (secondInsertVec[1]) begin // @[Sbuffer.scala 458:32]
        vtag_1 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_1 <= _GEN_287;
      end
    end else begin
      vtag_1 <= _GEN_287;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_2 <= _GEN_292;
      end else if (secondInsertVec[2]) begin // @[Sbuffer.scala 458:32]
        vtag_2 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_2 <= _GEN_292;
      end
    end else begin
      vtag_2 <= _GEN_292;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_3 <= _GEN_297;
      end else if (secondInsertVec[3]) begin // @[Sbuffer.scala 458:32]
        vtag_3 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_3 <= _GEN_297;
      end
    end else begin
      vtag_3 <= _GEN_297;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_4 <= _GEN_302;
      end else if (secondInsertVec[4]) begin // @[Sbuffer.scala 458:32]
        vtag_4 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_4 <= _GEN_302;
      end
    end else begin
      vtag_4 <= _GEN_302;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_5 <= _GEN_307;
      end else if (secondInsertVec[5]) begin // @[Sbuffer.scala 458:32]
        vtag_5 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_5 <= _GEN_307;
      end
    end else begin
      vtag_5 <= _GEN_307;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_6 <= _GEN_312;
      end else if (secondInsertVec[6]) begin // @[Sbuffer.scala 458:32]
        vtag_6 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_6 <= _GEN_312;
      end
    end else begin
      vtag_6 <= _GEN_312;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_7 <= _GEN_317;
      end else if (secondInsertVec[7]) begin // @[Sbuffer.scala 458:32]
        vtag_7 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_7 <= _GEN_317;
      end
    end else begin
      vtag_7 <= _GEN_317;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_8 <= _GEN_322;
      end else if (secondInsertVec[8]) begin // @[Sbuffer.scala 458:32]
        vtag_8 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_8 <= _GEN_322;
      end
    end else begin
      vtag_8 <= _GEN_322;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_9 <= _GEN_327;
      end else if (secondInsertVec[9]) begin // @[Sbuffer.scala 458:32]
        vtag_9 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_9 <= _GEN_327;
      end
    end else begin
      vtag_9 <= _GEN_327;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_10 <= _GEN_332;
      end else if (secondInsertVec[10]) begin // @[Sbuffer.scala 458:32]
        vtag_10 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_10 <= _GEN_332;
      end
    end else begin
      vtag_10 <= _GEN_332;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_11 <= _GEN_337;
      end else if (secondInsertVec[11]) begin // @[Sbuffer.scala 458:32]
        vtag_11 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_11 <= _GEN_337;
      end
    end else begin
      vtag_11 <= _GEN_337;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_12 <= _GEN_342;
      end else if (secondInsertVec[12]) begin // @[Sbuffer.scala 458:32]
        vtag_12 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_12 <= _GEN_342;
      end
    end else begin
      vtag_12 <= _GEN_342;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_13 <= _GEN_347;
      end else if (secondInsertVec[13]) begin // @[Sbuffer.scala 458:32]
        vtag_13 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_13 <= _GEN_347;
      end
    end else begin
      vtag_13 <= _GEN_347;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_14 <= _GEN_352;
      end else if (secondInsertVec[14]) begin // @[Sbuffer.scala 458:32]
        vtag_14 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_14 <= _GEN_352;
      end
    end else begin
      vtag_14 <= _GEN_352;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        vtag_15 <= _GEN_357;
      end else if (secondInsertVec[15]) begin // @[Sbuffer.scala 458:32]
        vtag_15 <= invtags_1; // @[Sbuffer.scala 467:24]
      end else begin
        vtag_15 <= _GEN_357;
      end
    end else begin
      vtag_15 <= _GEN_357;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_0 <= _GEN_280;
      end else if (secondInsertVec[0]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_0 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_0 <= _GEN_280;
        end
      end else begin
        waitInflightMask_0 <= _GEN_280;
      end
    end else begin
      waitInflightMask_0 <= _GEN_280;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_1 <= _GEN_285;
      end else if (secondInsertVec[1]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_1 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_1 <= _GEN_285;
        end
      end else begin
        waitInflightMask_1 <= _GEN_285;
      end
    end else begin
      waitInflightMask_1 <= _GEN_285;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_2 <= _GEN_290;
      end else if (secondInsertVec[2]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_2 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_2 <= _GEN_290;
        end
      end else begin
        waitInflightMask_2 <= _GEN_290;
      end
    end else begin
      waitInflightMask_2 <= _GEN_290;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_3 <= _GEN_295;
      end else if (secondInsertVec[3]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_3 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_3 <= _GEN_295;
        end
      end else begin
        waitInflightMask_3 <= _GEN_295;
      end
    end else begin
      waitInflightMask_3 <= _GEN_295;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_4 <= _GEN_300;
      end else if (secondInsertVec[4]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_4 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_4 <= _GEN_300;
        end
      end else begin
        waitInflightMask_4 <= _GEN_300;
      end
    end else begin
      waitInflightMask_4 <= _GEN_300;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_5 <= _GEN_305;
      end else if (secondInsertVec[5]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_5 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_5 <= _GEN_305;
        end
      end else begin
        waitInflightMask_5 <= _GEN_305;
      end
    end else begin
      waitInflightMask_5 <= _GEN_305;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_6 <= _GEN_310;
      end else if (secondInsertVec[6]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_6 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_6 <= _GEN_310;
        end
      end else begin
        waitInflightMask_6 <= _GEN_310;
      end
    end else begin
      waitInflightMask_6 <= _GEN_310;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_7 <= _GEN_315;
      end else if (secondInsertVec[7]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_7 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_7 <= _GEN_315;
        end
      end else begin
        waitInflightMask_7 <= _GEN_315;
      end
    end else begin
      waitInflightMask_7 <= _GEN_315;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_8 <= _GEN_320;
      end else if (secondInsertVec[8]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_8 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_8 <= _GEN_320;
        end
      end else begin
        waitInflightMask_8 <= _GEN_320;
      end
    end else begin
      waitInflightMask_8 <= _GEN_320;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_9 <= _GEN_325;
      end else if (secondInsertVec[9]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_9 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_9 <= _GEN_325;
        end
      end else begin
        waitInflightMask_9 <= _GEN_325;
      end
    end else begin
      waitInflightMask_9 <= _GEN_325;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_10 <= _GEN_330;
      end else if (secondInsertVec[10]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_10 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_10 <= _GEN_330;
        end
      end else begin
        waitInflightMask_10 <= _GEN_330;
      end
    end else begin
      waitInflightMask_10 <= _GEN_330;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_11 <= _GEN_335;
      end else if (secondInsertVec[11]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_11 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_11 <= _GEN_335;
        end
      end else begin
        waitInflightMask_11 <= _GEN_335;
      end
    end else begin
      waitInflightMask_11 <= _GEN_335;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_12 <= _GEN_340;
      end else if (secondInsertVec[12]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_12 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_12 <= _GEN_340;
        end
      end else begin
        waitInflightMask_12 <= _GEN_340;
      end
    end else begin
      waitInflightMask_12 <= _GEN_340;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_13 <= _GEN_345;
      end else if (secondInsertVec[13]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_13 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_13 <= _GEN_345;
        end
      end else begin
        waitInflightMask_13 <= _GEN_345;
      end
    end else begin
      waitInflightMask_13 <= _GEN_345;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_14 <= _GEN_350;
      end else if (secondInsertVec[14]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_14 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_14 <= _GEN_350;
        end
      end else begin
        waitInflightMask_14 <= _GEN_350;
      end
    end else begin
      waitInflightMask_14 <= _GEN_350;
    end
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        waitInflightMask_15 <= _GEN_355;
      end else if (secondInsertVec[15]) begin // @[Sbuffer.scala 458:32]
        if (_stateVec_0_w_sameblock_inflight_T_1) begin // @[Sbuffer.scala 461:40]
          waitInflightMask_15 <= sameBlockInflightMask_1; // @[Sbuffer.scala 462:38]
        end else begin
          waitInflightMask_15 <= _GEN_355;
        end
      end else begin
        waitInflightMask_15 <= _GEN_355;
      end
    end else begin
      waitInflightMask_15 <= _GEN_355;
    end
    missqReplayHasTimeOut_REG <= missqReplayTimeOutMask_0 | f_tail_27; // @[PriorityMuxDefault.scala 46:46]
    missqReplayHasTimeOut_REG_1 <= sbuffer_out_s0_valid & sbuffer_out_s0_cango; // @[Sbuffer.scala 652:47]
    if (missqReplayHasTimeOutGen) begin // @[Reg.scala 20:18]
      if (missqReplayTimeOutMask_0) begin // @[PriorityMuxDefault.scala 46:13]
        missqReplayTimeOutIdx <= 4'h0;
      end else if (missqReplayTimeOutMask_1) begin // @[PriorityMuxDefault.scala 46:13]
        missqReplayTimeOutIdx <= 4'h1;
      end else if (missqReplayTimeOutMask_2) begin // @[PriorityMuxDefault.scala 46:13]
        missqReplayTimeOutIdx <= 4'h2;
      end else begin
        missqReplayTimeOutIdx <= d_tail_25;
      end
    end
    do_uarch_drain_REG <= tag_mismatch_1 | tag_mismatch; // @[Sbuffer.scala 803:25 810:32]
    if (_dataModule_io_writeReq_1_valid_T) begin // @[Sbuffer.scala 511:20]
      if (canMerge_1) begin // @[Sbuffer.scala 512:24]
        if (mergeVec_1[15]) begin // @[Sbuffer.scala 482:32]
          do_uarch_drain_REG_1 <= _GEN_403;
        end else if (mergeVec_1[14]) begin // @[Sbuffer.scala 482:32]
          do_uarch_drain_REG_1 <= _GEN_400;
        end else begin
          do_uarch_drain_REG_1 <= _GEN_399;
        end
      end else begin
        do_uarch_drain_REG_1 <= _GEN_262;
      end
    end else begin
      do_uarch_drain_REG_1 <= _GEN_262;
    end
    do_uarch_drain_REG_2 <= do_uarch_drain_REG_1; // @[Sbuffer.scala 441:68]
    accessIdx_0_valid_REG <= io_in_0_ready & io_in_0_valid; // @[Decoupled.scala 51:35]
    if (canMerge_0) begin // @[Sbuffer.scala 510:37]
      if (mergeMask_0_0) begin // @[Mux.scala 47:70]
        accessIdx_0_bits_REG <= 4'h0;
      end else if (mergeMask_0_1) begin // @[Mux.scala 47:70]
        accessIdx_0_bits_REG <= 4'h1;
      end else if (mergeMask_0_2) begin // @[Mux.scala 47:70]
        accessIdx_0_bits_REG <= 4'h2;
      end else begin
        accessIdx_0_bits_REG <= _mergeIdx_T_11;
      end
    end else begin
      accessIdx_0_bits_REG <= insertIdx;
    end
    accessIdx_1_valid_REG <= io_in_1_ready & io_in_1_valid; // @[Decoupled.scala 51:35]
    if (canMerge_1) begin // @[Sbuffer.scala 510:37]
      if (mergeMask_1_0) begin // @[Mux.scala 47:70]
        accessIdx_1_bits_REG <= 4'h0;
      end else if (mergeMask_1_1) begin // @[Mux.scala 47:70]
        accessIdx_1_bits_REG <= 4'h1;
      end else if (mergeMask_1_2) begin // @[Mux.scala 47:70]
        accessIdx_1_bits_REG <= 4'h2;
      end else begin
        accessIdx_1_bits_REG <= _mergeIdx_T_25;
      end
    end else begin
      accessIdx_1_bits_REG <= insertIdx_1;
    end
    threshold <= io_csrCtrl_sbuffer_threshold + 4'h1; // @[Sbuffer.scala 549:56]
    io_flush_empty_REG <= empty & io_sqempty; // @[Sbuffer.scala 557:35]
    blockDcacheWrite <= |_shouldWaitWriteFinish_T_8; // @[Sbuffer.scala 662:13]
    if (sbuffer_out_s0_fire) begin // @[Reg.scala 20:18]
      if (missqReplayHasTimeOut) begin // @[Sbuffer.scala 634:39]
        sbuffer_out_s1_evictionIdx <= missqReplayTimeOutIdx;
      end else if (need_drain) begin // @[Sbuffer.scala 636:8]
        if (_candidateVec_T_1) begin // @[Mux.scala 47:70]
          sbuffer_out_s1_evictionIdx <= 4'h0;
        end else begin
          sbuffer_out_s1_evictionIdx <= _drainIdx_T_13;
        end
      end else if (cohHasTimeOut) begin // @[Sbuffer.scala 638:10]
        sbuffer_out_s1_evictionIdx <= cohTimeOutIdx;
      end else begin
        sbuffer_out_s1_evictionIdx <= Sbuffer_PLRU_io_replaceWay;
      end
    end
    if (sbuffer_out_s0_fire) begin // @[Reg.scala 20:18]
      if (4'hf == sbuffer_out_s0_evictionIdx) begin // @[Sbuffer.scala 595:53]
        sbuffer_out_s1_evictionPTag <= ptag_15; // @[Sbuffer.scala 595:53]
      end else if (4'he == sbuffer_out_s0_evictionIdx) begin // @[Sbuffer.scala 595:53]
        sbuffer_out_s1_evictionPTag <= ptag_14; // @[Sbuffer.scala 595:53]
      end else if (4'hd == sbuffer_out_s0_evictionIdx) begin // @[Sbuffer.scala 595:53]
        sbuffer_out_s1_evictionPTag <= ptag_13; // @[Sbuffer.scala 595:53]
      end else begin
        sbuffer_out_s1_evictionPTag <= _GEN_787;
      end
    end
    if (sbuffer_out_s0_fire) begin // @[Reg.scala 20:18]
      if (4'hf == sbuffer_out_s0_evictionIdx) begin // @[Reg.scala 20:22]
        sbuffer_out_s1_evictionVTag <= vtag_15; // @[Reg.scala 20:22]
      end else if (4'he == sbuffer_out_s0_evictionIdx) begin // @[Reg.scala 20:22]
        sbuffer_out_s1_evictionVTag <= vtag_14; // @[Reg.scala 20:22]
      end else if (4'hd == sbuffer_out_s0_evictionIdx) begin // @[Reg.scala 20:22]
        sbuffer_out_s1_evictionVTag <= vtag_13; // @[Reg.scala 20:22]
      end else begin
        sbuffer_out_s1_evictionVTag <= _GEN_903;
      end
    end
    REG <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_1 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_2 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_3 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_4 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_5 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_6 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_7 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_8 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_9 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_10 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_11 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_12 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_13 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_14 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_15 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_16 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_17 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_18 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_19 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_20 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_21 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_22 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_23 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_24 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_25 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_26 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_27 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_28 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_29 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_30 <= io_dcache_main_pipe_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_31 <= io_dcache_main_pipe_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_32 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_33 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_34 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_35 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_36 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_37 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_38 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_39 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_40 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_41 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_42 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_43 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_44 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_45 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_46 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_47 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_48 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_49 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_50 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_51 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_52 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_53 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_54 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_55 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_56 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_57 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_58 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_59 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_60 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_61 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    REG_62 <= io_dcache_refill_hit_resp_valid; // @[Sbuffer.scala 743:16]
    REG_63 <= io_dcache_refill_hit_resp_bits_id[3:0]; // @[Sbuffer.scala 720:7]
    tag_mismatch_REG <= io_forward_0_valid; // @[Sbuffer.scala 799:31]
    tag_mismatch_REG_31 <= vtag_15 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_30 <= ptag_15; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_31 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_32 <= _candidateVec_T_61 | stateVec_15_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_29 <= vtag_14 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_28 <= ptag_14; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_29 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_30 <= _candidateVec_T_57 | stateVec_14_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_27 <= vtag_13 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_26 <= ptag_13; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_27 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_28 <= _candidateVec_T_53 | stateVec_13_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_25 <= vtag_12 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_24 <= ptag_12; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_25 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_26 <= _candidateVec_T_49 | stateVec_12_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_23 <= vtag_11 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_22 <= ptag_11; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_23 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_24 <= _candidateVec_T_45 | stateVec_11_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_21 <= vtag_10 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_20 <= ptag_10; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_21 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_22 <= _candidateVec_T_41 | stateVec_10_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_19 <= vtag_9 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_18 <= ptag_9; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_19 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_20 <= _candidateVec_T_37 | stateVec_9_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_17 <= vtag_8 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_16 <= ptag_8; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_17 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_18 <= _candidateVec_T_33 | stateVec_8_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_15 <= vtag_7 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_14 <= ptag_7; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_15 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_16 <= _candidateVec_T_29 | stateVec_7_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_13 <= vtag_6 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_12 <= ptag_6; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_13 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_14 <= _candidateVec_T_25 | stateVec_6_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_11 <= vtag_5 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_10 <= ptag_5; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_11 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_12 <= _candidateVec_T_21 | stateVec_5_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_9 <= vtag_4 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_8 <= ptag_4; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_9 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_10 <= _candidateVec_T_17 | stateVec_4_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_7 <= vtag_3 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_6 <= ptag_3; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_7 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_8 <= _candidateVec_T_13 | stateVec_3_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_5 <= vtag_2 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_4 <= ptag_2; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_5 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_6 <= _candidateVec_T_9 | stateVec_2_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_3 <= vtag_1 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_2 <= ptag_1; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_3 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_4 <= _candidateVec_T_5 | stateVec_1_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_1 <= vtag_0 == io_forward_0_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r <= ptag_0; // @[Reg.scala 20:22]
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_1 <= io_forward_0_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_2 <= _candidateVec_T_1 | stateVec_0_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_33 <= io_forward_1_valid; // @[Sbuffer.scala 799:31]
    tag_mismatch_REG_64 <= vtag_15 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_62 <= ptag_15; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_63 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_65 <= _candidateVec_T_61 | stateVec_15_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_62 <= vtag_14 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_60 <= ptag_14; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_61 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_63 <= _candidateVec_T_57 | stateVec_14_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_60 <= vtag_13 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_58 <= ptag_13; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_59 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_61 <= _candidateVec_T_53 | stateVec_13_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_58 <= vtag_12 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_56 <= ptag_12; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_57 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_59 <= _candidateVec_T_49 | stateVec_12_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_56 <= vtag_11 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_54 <= ptag_11; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_55 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_57 <= _candidateVec_T_45 | stateVec_11_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_54 <= vtag_10 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_52 <= ptag_10; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_53 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_55 <= _candidateVec_T_41 | stateVec_10_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_52 <= vtag_9 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_50 <= ptag_9; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_51 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_53 <= _candidateVec_T_37 | stateVec_9_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_50 <= vtag_8 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_48 <= ptag_8; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_49 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_51 <= _candidateVec_T_33 | stateVec_8_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_48 <= vtag_7 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_46 <= ptag_7; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_47 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_49 <= _candidateVec_T_29 | stateVec_7_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_46 <= vtag_6 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_44 <= ptag_6; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_45 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_47 <= _candidateVec_T_25 | stateVec_6_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_44 <= vtag_5 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_42 <= ptag_5; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_43 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_45 <= _candidateVec_T_21 | stateVec_5_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_42 <= vtag_4 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_40 <= ptag_4; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_41 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_43 <= _candidateVec_T_17 | stateVec_4_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_40 <= vtag_3 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_38 <= ptag_3; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_39 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_41 <= _candidateVec_T_13 | stateVec_3_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_38 <= vtag_2 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_36 <= ptag_2; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_37 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_39 <= _candidateVec_T_9 | stateVec_2_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_36 <= vtag_1 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_34 <= ptag_1; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_35 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_37 <= _candidateVec_T_5 | stateVec_1_state_inflight; // @[Sbuffer.scala 800:78]
    tag_mismatch_REG_34 <= vtag_0 == io_forward_1_vaddr[38:6]; // @[Sbuffer.scala 795:54]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_32 <= ptag_0; // @[Reg.scala 20:22]
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      ptag_matches_r_33 <= io_forward_1_paddr[35:6]; // @[Reg.scala 20:22]
    end
    tag_mismatch_REG_35 <= _candidateVec_T_1 | stateVec_0_state_inflight; // @[Sbuffer.scala 800:78]
    valid_tag_match_reg_0 <= vtag_matches__0 & _candidateVec_T_1; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_1 <= vtag_matches__1 & _candidateVec_T_5; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_2 <= vtag_matches__2 & _candidateVec_T_9; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_3 <= vtag_matches__3 & _candidateVec_T_13; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_4 <= vtag_matches__4 & _candidateVec_T_17; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_5 <= vtag_matches__5 & _candidateVec_T_21; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_6 <= vtag_matches__6 & _candidateVec_T_25; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_7 <= vtag_matches__7 & _candidateVec_T_29; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_8 <= vtag_matches__8 & _candidateVec_T_33; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_9 <= vtag_matches__9 & _candidateVec_T_37; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_10 <= vtag_matches__10 & _candidateVec_T_41; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_11 <= vtag_matches__11 & _candidateVec_T_45; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_12 <= vtag_matches__12 & _candidateVec_T_49; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_13 <= vtag_matches__13 & _candidateVec_T_53; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_14 <= vtag_matches__14 & _candidateVec_T_57; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_15 <= vtag_matches__15 & _candidateVec_T_61; // @[Sbuffer.scala 812:58]
    inflight_tag_match_reg_0 <= vtag_matches__0 & stateVec_0_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_1 <= vtag_matches__1 & stateVec_1_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_2 <= vtag_matches__2 & stateVec_2_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_3 <= vtag_matches__3 & stateVec_3_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_4 <= vtag_matches__4 & stateVec_4_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_5 <= vtag_matches__5 & stateVec_5_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_6 <= vtag_matches__6 & stateVec_6_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_7 <= vtag_matches__7 & stateVec_7_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_8 <= vtag_matches__8 & stateVec_8_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_9 <= vtag_matches__9 & stateVec_9_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_10 <= vtag_matches__10 & stateVec_10_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_11 <= vtag_matches__11 & stateVec_11_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_12 <= vtag_matches__12 & stateVec_12_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_13 <= vtag_matches__13 & stateVec_13_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_14 <= vtag_matches__14 & stateVec_14_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_15 <= vtag_matches__15 & stateVec_15_state_inflight; // @[Sbuffer.scala 813:61]
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_0 <= dataModule_io_maskOut_0_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_0 <= dataModule_io_maskOut_0_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_0 <= dataModule_io_maskOut_0_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_0 <= _GEN_3297;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_1 <= dataModule_io_maskOut_0_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_1 <= dataModule_io_maskOut_0_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_1 <= dataModule_io_maskOut_0_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_1 <= _GEN_3305;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_2 <= dataModule_io_maskOut_0_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_2 <= dataModule_io_maskOut_0_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_2 <= dataModule_io_maskOut_0_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_2 <= _GEN_3313;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_3 <= dataModule_io_maskOut_0_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_3 <= dataModule_io_maskOut_0_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_3 <= dataModule_io_maskOut_0_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_3 <= _GEN_3321;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_4 <= dataModule_io_maskOut_0_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_4 <= dataModule_io_maskOut_0_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_4 <= dataModule_io_maskOut_0_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_4 <= _GEN_3329;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_5 <= dataModule_io_maskOut_0_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_5 <= dataModule_io_maskOut_0_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_5 <= dataModule_io_maskOut_0_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_5 <= _GEN_3337;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_6 <= dataModule_io_maskOut_0_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_6 <= dataModule_io_maskOut_0_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_6 <= dataModule_io_maskOut_0_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_6 <= _GEN_3345;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_7 <= dataModule_io_maskOut_0_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_7 <= dataModule_io_maskOut_0_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__0_7 <= dataModule_io_maskOut_0_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__0_7 <= _GEN_3353;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_0 <= dataModule_io_maskOut_1_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_0 <= dataModule_io_maskOut_1_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_0 <= dataModule_io_maskOut_1_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_0 <= _GEN_3361;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_1 <= dataModule_io_maskOut_1_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_1 <= dataModule_io_maskOut_1_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_1 <= dataModule_io_maskOut_1_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_1 <= _GEN_3369;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_2 <= dataModule_io_maskOut_1_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_2 <= dataModule_io_maskOut_1_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_2 <= dataModule_io_maskOut_1_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_2 <= _GEN_3377;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_3 <= dataModule_io_maskOut_1_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_3 <= dataModule_io_maskOut_1_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_3 <= dataModule_io_maskOut_1_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_3 <= _GEN_3385;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_4 <= dataModule_io_maskOut_1_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_4 <= dataModule_io_maskOut_1_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_4 <= dataModule_io_maskOut_1_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_4 <= _GEN_3393;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_5 <= dataModule_io_maskOut_1_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_5 <= dataModule_io_maskOut_1_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_5 <= dataModule_io_maskOut_1_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_5 <= _GEN_3401;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_6 <= dataModule_io_maskOut_1_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_6 <= dataModule_io_maskOut_1_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_6 <= dataModule_io_maskOut_1_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_6 <= _GEN_3409;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_7 <= dataModule_io_maskOut_1_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_7 <= dataModule_io_maskOut_1_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__1_7 <= dataModule_io_maskOut_1_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__1_7 <= _GEN_3417;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_0 <= dataModule_io_maskOut_2_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_0 <= dataModule_io_maskOut_2_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_0 <= dataModule_io_maskOut_2_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_0 <= _GEN_3425;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_1 <= dataModule_io_maskOut_2_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_1 <= dataModule_io_maskOut_2_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_1 <= dataModule_io_maskOut_2_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_1 <= _GEN_3433;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_2 <= dataModule_io_maskOut_2_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_2 <= dataModule_io_maskOut_2_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_2 <= dataModule_io_maskOut_2_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_2 <= _GEN_3441;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_3 <= dataModule_io_maskOut_2_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_3 <= dataModule_io_maskOut_2_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_3 <= dataModule_io_maskOut_2_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_3 <= _GEN_3449;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_4 <= dataModule_io_maskOut_2_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_4 <= dataModule_io_maskOut_2_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_4 <= dataModule_io_maskOut_2_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_4 <= _GEN_3457;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_5 <= dataModule_io_maskOut_2_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_5 <= dataModule_io_maskOut_2_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_5 <= dataModule_io_maskOut_2_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_5 <= _GEN_3465;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_6 <= dataModule_io_maskOut_2_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_6 <= dataModule_io_maskOut_2_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_6 <= dataModule_io_maskOut_2_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_6 <= _GEN_3473;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_7 <= dataModule_io_maskOut_2_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_7 <= dataModule_io_maskOut_2_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__2_7 <= dataModule_io_maskOut_2_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__2_7 <= _GEN_3481;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_0 <= dataModule_io_maskOut_3_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_0 <= dataModule_io_maskOut_3_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_0 <= dataModule_io_maskOut_3_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_0 <= _GEN_3489;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_1 <= dataModule_io_maskOut_3_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_1 <= dataModule_io_maskOut_3_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_1 <= dataModule_io_maskOut_3_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_1 <= _GEN_3497;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_2 <= dataModule_io_maskOut_3_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_2 <= dataModule_io_maskOut_3_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_2 <= dataModule_io_maskOut_3_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_2 <= _GEN_3505;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_3 <= dataModule_io_maskOut_3_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_3 <= dataModule_io_maskOut_3_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_3 <= dataModule_io_maskOut_3_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_3 <= _GEN_3513;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_4 <= dataModule_io_maskOut_3_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_4 <= dataModule_io_maskOut_3_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_4 <= dataModule_io_maskOut_3_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_4 <= _GEN_3521;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_5 <= dataModule_io_maskOut_3_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_5 <= dataModule_io_maskOut_3_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_5 <= dataModule_io_maskOut_3_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_5 <= _GEN_3529;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_6 <= dataModule_io_maskOut_3_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_6 <= dataModule_io_maskOut_3_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_6 <= dataModule_io_maskOut_3_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_6 <= _GEN_3537;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_7 <= dataModule_io_maskOut_3_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_7 <= dataModule_io_maskOut_3_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__3_7 <= dataModule_io_maskOut_3_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__3_7 <= _GEN_3545;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_0 <= dataModule_io_maskOut_4_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_0 <= dataModule_io_maskOut_4_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_0 <= dataModule_io_maskOut_4_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_0 <= _GEN_3553;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_1 <= dataModule_io_maskOut_4_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_1 <= dataModule_io_maskOut_4_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_1 <= dataModule_io_maskOut_4_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_1 <= _GEN_3561;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_2 <= dataModule_io_maskOut_4_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_2 <= dataModule_io_maskOut_4_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_2 <= dataModule_io_maskOut_4_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_2 <= _GEN_3569;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_3 <= dataModule_io_maskOut_4_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_3 <= dataModule_io_maskOut_4_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_3 <= dataModule_io_maskOut_4_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_3 <= _GEN_3577;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_4 <= dataModule_io_maskOut_4_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_4 <= dataModule_io_maskOut_4_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_4 <= dataModule_io_maskOut_4_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_4 <= _GEN_3585;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_5 <= dataModule_io_maskOut_4_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_5 <= dataModule_io_maskOut_4_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_5 <= dataModule_io_maskOut_4_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_5 <= _GEN_3593;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_6 <= dataModule_io_maskOut_4_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_6 <= dataModule_io_maskOut_4_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_6 <= dataModule_io_maskOut_4_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_6 <= _GEN_3601;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_7 <= dataModule_io_maskOut_4_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_7 <= dataModule_io_maskOut_4_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__4_7 <= dataModule_io_maskOut_4_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__4_7 <= _GEN_3609;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_0 <= dataModule_io_maskOut_5_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_0 <= dataModule_io_maskOut_5_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_0 <= dataModule_io_maskOut_5_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_0 <= _GEN_3617;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_1 <= dataModule_io_maskOut_5_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_1 <= dataModule_io_maskOut_5_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_1 <= dataModule_io_maskOut_5_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_1 <= _GEN_3625;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_2 <= dataModule_io_maskOut_5_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_2 <= dataModule_io_maskOut_5_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_2 <= dataModule_io_maskOut_5_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_2 <= _GEN_3633;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_3 <= dataModule_io_maskOut_5_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_3 <= dataModule_io_maskOut_5_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_3 <= dataModule_io_maskOut_5_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_3 <= _GEN_3641;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_4 <= dataModule_io_maskOut_5_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_4 <= dataModule_io_maskOut_5_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_4 <= dataModule_io_maskOut_5_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_4 <= _GEN_3649;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_5 <= dataModule_io_maskOut_5_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_5 <= dataModule_io_maskOut_5_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_5 <= dataModule_io_maskOut_5_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_5 <= _GEN_3657;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_6 <= dataModule_io_maskOut_5_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_6 <= dataModule_io_maskOut_5_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_6 <= dataModule_io_maskOut_5_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_6 <= _GEN_3665;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_7 <= dataModule_io_maskOut_5_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_7 <= dataModule_io_maskOut_5_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__5_7 <= dataModule_io_maskOut_5_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__5_7 <= _GEN_3673;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_0 <= dataModule_io_maskOut_6_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_0 <= dataModule_io_maskOut_6_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_0 <= dataModule_io_maskOut_6_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_0 <= _GEN_3681;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_1 <= dataModule_io_maskOut_6_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_1 <= dataModule_io_maskOut_6_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_1 <= dataModule_io_maskOut_6_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_1 <= _GEN_3689;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_2 <= dataModule_io_maskOut_6_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_2 <= dataModule_io_maskOut_6_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_2 <= dataModule_io_maskOut_6_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_2 <= _GEN_3697;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_3 <= dataModule_io_maskOut_6_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_3 <= dataModule_io_maskOut_6_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_3 <= dataModule_io_maskOut_6_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_3 <= _GEN_3705;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_4 <= dataModule_io_maskOut_6_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_4 <= dataModule_io_maskOut_6_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_4 <= dataModule_io_maskOut_6_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_4 <= _GEN_3713;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_5 <= dataModule_io_maskOut_6_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_5 <= dataModule_io_maskOut_6_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_5 <= dataModule_io_maskOut_6_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_5 <= _GEN_3721;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_6 <= dataModule_io_maskOut_6_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_6 <= dataModule_io_maskOut_6_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_6 <= dataModule_io_maskOut_6_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_6 <= _GEN_3729;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_7 <= dataModule_io_maskOut_6_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_7 <= dataModule_io_maskOut_6_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__6_7 <= dataModule_io_maskOut_6_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__6_7 <= _GEN_3737;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_0 <= dataModule_io_maskOut_7_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_0 <= dataModule_io_maskOut_7_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_0 <= dataModule_io_maskOut_7_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_0 <= _GEN_3745;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_1 <= dataModule_io_maskOut_7_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_1 <= dataModule_io_maskOut_7_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_1 <= dataModule_io_maskOut_7_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_1 <= _GEN_3753;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_2 <= dataModule_io_maskOut_7_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_2 <= dataModule_io_maskOut_7_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_2 <= dataModule_io_maskOut_7_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_2 <= _GEN_3761;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_3 <= dataModule_io_maskOut_7_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_3 <= dataModule_io_maskOut_7_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_3 <= dataModule_io_maskOut_7_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_3 <= _GEN_3769;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_4 <= dataModule_io_maskOut_7_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_4 <= dataModule_io_maskOut_7_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_4 <= dataModule_io_maskOut_7_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_4 <= _GEN_3777;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_5 <= dataModule_io_maskOut_7_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_5 <= dataModule_io_maskOut_7_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_5 <= dataModule_io_maskOut_7_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_5 <= _GEN_3785;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_6 <= dataModule_io_maskOut_7_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_6 <= dataModule_io_maskOut_7_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_6 <= dataModule_io_maskOut_7_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_6 <= _GEN_3793;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_7 <= dataModule_io_maskOut_7_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_7 <= dataModule_io_maskOut_7_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__7_7 <= dataModule_io_maskOut_7_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__7_7 <= _GEN_3801;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_0 <= dataModule_io_maskOut_8_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_0 <= dataModule_io_maskOut_8_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_0 <= dataModule_io_maskOut_8_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_0 <= _GEN_3809;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_1 <= dataModule_io_maskOut_8_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_1 <= dataModule_io_maskOut_8_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_1 <= dataModule_io_maskOut_8_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_1 <= _GEN_3817;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_2 <= dataModule_io_maskOut_8_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_2 <= dataModule_io_maskOut_8_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_2 <= dataModule_io_maskOut_8_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_2 <= _GEN_3825;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_3 <= dataModule_io_maskOut_8_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_3 <= dataModule_io_maskOut_8_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_3 <= dataModule_io_maskOut_8_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_3 <= _GEN_3833;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_4 <= dataModule_io_maskOut_8_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_4 <= dataModule_io_maskOut_8_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_4 <= dataModule_io_maskOut_8_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_4 <= _GEN_3841;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_5 <= dataModule_io_maskOut_8_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_5 <= dataModule_io_maskOut_8_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_5 <= dataModule_io_maskOut_8_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_5 <= _GEN_3849;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_6 <= dataModule_io_maskOut_8_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_6 <= dataModule_io_maskOut_8_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_6 <= dataModule_io_maskOut_8_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_6 <= _GEN_3857;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_7 <= dataModule_io_maskOut_8_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_7 <= dataModule_io_maskOut_8_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__8_7 <= dataModule_io_maskOut_8_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__8_7 <= _GEN_3865;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_0 <= dataModule_io_maskOut_9_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_0 <= dataModule_io_maskOut_9_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_0 <= dataModule_io_maskOut_9_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_0 <= _GEN_3873;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_1 <= dataModule_io_maskOut_9_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_1 <= dataModule_io_maskOut_9_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_1 <= dataModule_io_maskOut_9_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_1 <= _GEN_3881;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_2 <= dataModule_io_maskOut_9_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_2 <= dataModule_io_maskOut_9_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_2 <= dataModule_io_maskOut_9_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_2 <= _GEN_3889;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_3 <= dataModule_io_maskOut_9_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_3 <= dataModule_io_maskOut_9_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_3 <= dataModule_io_maskOut_9_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_3 <= _GEN_3897;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_4 <= dataModule_io_maskOut_9_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_4 <= dataModule_io_maskOut_9_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_4 <= dataModule_io_maskOut_9_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_4 <= _GEN_3905;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_5 <= dataModule_io_maskOut_9_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_5 <= dataModule_io_maskOut_9_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_5 <= dataModule_io_maskOut_9_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_5 <= _GEN_3913;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_6 <= dataModule_io_maskOut_9_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_6 <= dataModule_io_maskOut_9_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_6 <= dataModule_io_maskOut_9_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_6 <= _GEN_3921;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_7 <= dataModule_io_maskOut_9_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_7 <= dataModule_io_maskOut_9_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__9_7 <= dataModule_io_maskOut_9_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__9_7 <= _GEN_3929;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_0 <= dataModule_io_maskOut_10_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_0 <= dataModule_io_maskOut_10_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_0 <= dataModule_io_maskOut_10_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_0 <= _GEN_3937;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_1 <= dataModule_io_maskOut_10_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_1 <= dataModule_io_maskOut_10_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_1 <= dataModule_io_maskOut_10_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_1 <= _GEN_3945;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_2 <= dataModule_io_maskOut_10_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_2 <= dataModule_io_maskOut_10_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_2 <= dataModule_io_maskOut_10_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_2 <= _GEN_3953;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_3 <= dataModule_io_maskOut_10_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_3 <= dataModule_io_maskOut_10_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_3 <= dataModule_io_maskOut_10_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_3 <= _GEN_3961;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_4 <= dataModule_io_maskOut_10_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_4 <= dataModule_io_maskOut_10_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_4 <= dataModule_io_maskOut_10_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_4 <= _GEN_3969;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_5 <= dataModule_io_maskOut_10_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_5 <= dataModule_io_maskOut_10_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_5 <= dataModule_io_maskOut_10_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_5 <= _GEN_3977;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_6 <= dataModule_io_maskOut_10_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_6 <= dataModule_io_maskOut_10_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_6 <= dataModule_io_maskOut_10_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_6 <= _GEN_3985;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_7 <= dataModule_io_maskOut_10_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_7 <= dataModule_io_maskOut_10_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__10_7 <= dataModule_io_maskOut_10_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__10_7 <= _GEN_3993;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_0 <= dataModule_io_maskOut_11_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_0 <= dataModule_io_maskOut_11_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_0 <= dataModule_io_maskOut_11_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_0 <= _GEN_4001;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_1 <= dataModule_io_maskOut_11_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_1 <= dataModule_io_maskOut_11_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_1 <= dataModule_io_maskOut_11_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_1 <= _GEN_4009;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_2 <= dataModule_io_maskOut_11_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_2 <= dataModule_io_maskOut_11_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_2 <= dataModule_io_maskOut_11_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_2 <= _GEN_4017;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_3 <= dataModule_io_maskOut_11_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_3 <= dataModule_io_maskOut_11_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_3 <= dataModule_io_maskOut_11_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_3 <= _GEN_4025;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_4 <= dataModule_io_maskOut_11_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_4 <= dataModule_io_maskOut_11_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_4 <= dataModule_io_maskOut_11_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_4 <= _GEN_4033;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_5 <= dataModule_io_maskOut_11_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_5 <= dataModule_io_maskOut_11_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_5 <= dataModule_io_maskOut_11_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_5 <= _GEN_4041;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_6 <= dataModule_io_maskOut_11_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_6 <= dataModule_io_maskOut_11_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_6 <= dataModule_io_maskOut_11_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_6 <= _GEN_4049;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_7 <= dataModule_io_maskOut_11_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_7 <= dataModule_io_maskOut_11_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__11_7 <= dataModule_io_maskOut_11_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__11_7 <= _GEN_4057;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_0 <= dataModule_io_maskOut_12_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_0 <= dataModule_io_maskOut_12_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_0 <= dataModule_io_maskOut_12_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_0 <= _GEN_4065;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_1 <= dataModule_io_maskOut_12_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_1 <= dataModule_io_maskOut_12_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_1 <= dataModule_io_maskOut_12_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_1 <= _GEN_4073;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_2 <= dataModule_io_maskOut_12_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_2 <= dataModule_io_maskOut_12_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_2 <= dataModule_io_maskOut_12_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_2 <= _GEN_4081;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_3 <= dataModule_io_maskOut_12_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_3 <= dataModule_io_maskOut_12_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_3 <= dataModule_io_maskOut_12_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_3 <= _GEN_4089;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_4 <= dataModule_io_maskOut_12_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_4 <= dataModule_io_maskOut_12_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_4 <= dataModule_io_maskOut_12_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_4 <= _GEN_4097;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_5 <= dataModule_io_maskOut_12_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_5 <= dataModule_io_maskOut_12_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_5 <= dataModule_io_maskOut_12_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_5 <= _GEN_4105;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_6 <= dataModule_io_maskOut_12_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_6 <= dataModule_io_maskOut_12_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_6 <= dataModule_io_maskOut_12_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_6 <= _GEN_4113;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_7 <= dataModule_io_maskOut_12_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_7 <= dataModule_io_maskOut_12_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__12_7 <= dataModule_io_maskOut_12_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__12_7 <= _GEN_4121;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_0 <= dataModule_io_maskOut_13_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_0 <= dataModule_io_maskOut_13_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_0 <= dataModule_io_maskOut_13_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_0 <= _GEN_4129;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_1 <= dataModule_io_maskOut_13_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_1 <= dataModule_io_maskOut_13_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_1 <= dataModule_io_maskOut_13_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_1 <= _GEN_4137;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_2 <= dataModule_io_maskOut_13_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_2 <= dataModule_io_maskOut_13_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_2 <= dataModule_io_maskOut_13_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_2 <= _GEN_4145;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_3 <= dataModule_io_maskOut_13_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_3 <= dataModule_io_maskOut_13_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_3 <= dataModule_io_maskOut_13_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_3 <= _GEN_4153;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_4 <= dataModule_io_maskOut_13_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_4 <= dataModule_io_maskOut_13_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_4 <= dataModule_io_maskOut_13_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_4 <= _GEN_4161;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_5 <= dataModule_io_maskOut_13_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_5 <= dataModule_io_maskOut_13_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_5 <= dataModule_io_maskOut_13_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_5 <= _GEN_4169;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_6 <= dataModule_io_maskOut_13_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_6 <= dataModule_io_maskOut_13_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_6 <= dataModule_io_maskOut_13_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_6 <= _GEN_4177;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_7 <= dataModule_io_maskOut_13_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_7 <= dataModule_io_maskOut_13_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__13_7 <= dataModule_io_maskOut_13_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__13_7 <= _GEN_4185;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_0 <= dataModule_io_maskOut_14_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_0 <= dataModule_io_maskOut_14_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_0 <= dataModule_io_maskOut_14_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_0 <= _GEN_4193;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_1 <= dataModule_io_maskOut_14_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_1 <= dataModule_io_maskOut_14_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_1 <= dataModule_io_maskOut_14_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_1 <= _GEN_4201;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_2 <= dataModule_io_maskOut_14_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_2 <= dataModule_io_maskOut_14_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_2 <= dataModule_io_maskOut_14_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_2 <= _GEN_4209;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_3 <= dataModule_io_maskOut_14_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_3 <= dataModule_io_maskOut_14_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_3 <= dataModule_io_maskOut_14_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_3 <= _GEN_4217;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_4 <= dataModule_io_maskOut_14_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_4 <= dataModule_io_maskOut_14_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_4 <= dataModule_io_maskOut_14_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_4 <= _GEN_4225;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_5 <= dataModule_io_maskOut_14_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_5 <= dataModule_io_maskOut_14_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_5 <= dataModule_io_maskOut_14_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_5 <= _GEN_4233;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_6 <= dataModule_io_maskOut_14_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_6 <= dataModule_io_maskOut_14_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_6 <= dataModule_io_maskOut_14_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_6 <= _GEN_4241;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_7 <= dataModule_io_maskOut_14_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_7 <= dataModule_io_maskOut_14_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__14_7 <= dataModule_io_maskOut_14_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__14_7 <= _GEN_4249;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_0 <= dataModule_io_maskOut_15_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_0 <= dataModule_io_maskOut_15_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_0 <= dataModule_io_maskOut_15_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_0 <= _GEN_4257;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_1 <= dataModule_io_maskOut_15_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_1 <= dataModule_io_maskOut_15_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_1 <= dataModule_io_maskOut_15_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_1 <= _GEN_4265;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_2 <= dataModule_io_maskOut_15_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_2 <= dataModule_io_maskOut_15_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_2 <= dataModule_io_maskOut_15_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_2 <= _GEN_4273;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_3 <= dataModule_io_maskOut_15_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_3 <= dataModule_io_maskOut_15_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_3 <= dataModule_io_maskOut_15_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_3 <= _GEN_4281;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_4 <= dataModule_io_maskOut_15_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_4 <= dataModule_io_maskOut_15_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_4 <= dataModule_io_maskOut_15_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_4 <= _GEN_4289;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_5 <= dataModule_io_maskOut_15_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_5 <= dataModule_io_maskOut_15_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_5 <= dataModule_io_maskOut_15_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_5 <= _GEN_4297;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_6 <= dataModule_io_maskOut_15_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_6 <= dataModule_io_maskOut_15_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_6 <= dataModule_io_maskOut_15_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_6 <= _GEN_4305;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_7 <= dataModule_io_maskOut_15_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_7 <= dataModule_io_maskOut_15_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg__15_7 <= dataModule_io_maskOut_15_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg__15_7 <= _GEN_4313;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_0 <= dataModule_io_dataOut_0_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_0 <= dataModule_io_dataOut_0_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_0 <= dataModule_io_dataOut_0_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_0 <= _GEN_4449;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_1 <= dataModule_io_dataOut_0_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_1 <= dataModule_io_dataOut_0_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_1 <= dataModule_io_dataOut_0_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_1 <= _GEN_4457;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_2 <= dataModule_io_dataOut_0_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_2 <= dataModule_io_dataOut_0_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_2 <= dataModule_io_dataOut_0_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_2 <= _GEN_4465;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_3 <= dataModule_io_dataOut_0_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_3 <= dataModule_io_dataOut_0_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_3 <= dataModule_io_dataOut_0_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_3 <= _GEN_4473;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_4 <= dataModule_io_dataOut_0_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_4 <= dataModule_io_dataOut_0_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_4 <= dataModule_io_dataOut_0_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_4 <= _GEN_4481;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_5 <= dataModule_io_dataOut_0_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_5 <= dataModule_io_dataOut_0_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_5 <= dataModule_io_dataOut_0_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_5 <= _GEN_4489;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_6 <= dataModule_io_dataOut_0_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_6 <= dataModule_io_dataOut_0_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_6 <= dataModule_io_dataOut_0_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_6 <= _GEN_4497;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_7 <= dataModule_io_dataOut_0_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_7 <= dataModule_io_dataOut_0_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__0_7 <= dataModule_io_dataOut_0_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__0_7 <= _GEN_4505;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_0 <= dataModule_io_dataOut_1_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_0 <= dataModule_io_dataOut_1_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_0 <= dataModule_io_dataOut_1_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_0 <= _GEN_4513;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_1 <= dataModule_io_dataOut_1_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_1 <= dataModule_io_dataOut_1_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_1 <= dataModule_io_dataOut_1_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_1 <= _GEN_4521;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_2 <= dataModule_io_dataOut_1_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_2 <= dataModule_io_dataOut_1_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_2 <= dataModule_io_dataOut_1_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_2 <= _GEN_4529;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_3 <= dataModule_io_dataOut_1_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_3 <= dataModule_io_dataOut_1_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_3 <= dataModule_io_dataOut_1_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_3 <= _GEN_4537;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_4 <= dataModule_io_dataOut_1_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_4 <= dataModule_io_dataOut_1_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_4 <= dataModule_io_dataOut_1_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_4 <= _GEN_4545;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_5 <= dataModule_io_dataOut_1_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_5 <= dataModule_io_dataOut_1_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_5 <= dataModule_io_dataOut_1_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_5 <= _GEN_4553;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_6 <= dataModule_io_dataOut_1_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_6 <= dataModule_io_dataOut_1_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_6 <= dataModule_io_dataOut_1_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_6 <= _GEN_4561;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_7 <= dataModule_io_dataOut_1_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_7 <= dataModule_io_dataOut_1_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__1_7 <= dataModule_io_dataOut_1_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__1_7 <= _GEN_4569;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_0 <= dataModule_io_dataOut_2_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_0 <= dataModule_io_dataOut_2_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_0 <= dataModule_io_dataOut_2_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_0 <= _GEN_4577;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_1 <= dataModule_io_dataOut_2_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_1 <= dataModule_io_dataOut_2_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_1 <= dataModule_io_dataOut_2_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_1 <= _GEN_4585;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_2 <= dataModule_io_dataOut_2_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_2 <= dataModule_io_dataOut_2_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_2 <= dataModule_io_dataOut_2_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_2 <= _GEN_4593;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_3 <= dataModule_io_dataOut_2_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_3 <= dataModule_io_dataOut_2_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_3 <= dataModule_io_dataOut_2_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_3 <= _GEN_4601;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_4 <= dataModule_io_dataOut_2_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_4 <= dataModule_io_dataOut_2_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_4 <= dataModule_io_dataOut_2_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_4 <= _GEN_4609;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_5 <= dataModule_io_dataOut_2_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_5 <= dataModule_io_dataOut_2_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_5 <= dataModule_io_dataOut_2_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_5 <= _GEN_4617;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_6 <= dataModule_io_dataOut_2_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_6 <= dataModule_io_dataOut_2_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_6 <= dataModule_io_dataOut_2_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_6 <= _GEN_4625;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_7 <= dataModule_io_dataOut_2_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_7 <= dataModule_io_dataOut_2_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__2_7 <= dataModule_io_dataOut_2_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__2_7 <= _GEN_4633;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_0 <= dataModule_io_dataOut_3_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_0 <= dataModule_io_dataOut_3_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_0 <= dataModule_io_dataOut_3_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_0 <= _GEN_4641;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_1 <= dataModule_io_dataOut_3_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_1 <= dataModule_io_dataOut_3_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_1 <= dataModule_io_dataOut_3_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_1 <= _GEN_4649;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_2 <= dataModule_io_dataOut_3_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_2 <= dataModule_io_dataOut_3_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_2 <= dataModule_io_dataOut_3_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_2 <= _GEN_4657;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_3 <= dataModule_io_dataOut_3_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_3 <= dataModule_io_dataOut_3_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_3 <= dataModule_io_dataOut_3_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_3 <= _GEN_4665;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_4 <= dataModule_io_dataOut_3_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_4 <= dataModule_io_dataOut_3_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_4 <= dataModule_io_dataOut_3_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_4 <= _GEN_4673;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_5 <= dataModule_io_dataOut_3_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_5 <= dataModule_io_dataOut_3_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_5 <= dataModule_io_dataOut_3_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_5 <= _GEN_4681;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_6 <= dataModule_io_dataOut_3_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_6 <= dataModule_io_dataOut_3_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_6 <= dataModule_io_dataOut_3_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_6 <= _GEN_4689;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_7 <= dataModule_io_dataOut_3_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_7 <= dataModule_io_dataOut_3_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__3_7 <= dataModule_io_dataOut_3_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__3_7 <= _GEN_4697;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_0 <= dataModule_io_dataOut_4_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_0 <= dataModule_io_dataOut_4_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_0 <= dataModule_io_dataOut_4_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_0 <= _GEN_4705;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_1 <= dataModule_io_dataOut_4_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_1 <= dataModule_io_dataOut_4_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_1 <= dataModule_io_dataOut_4_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_1 <= _GEN_4713;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_2 <= dataModule_io_dataOut_4_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_2 <= dataModule_io_dataOut_4_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_2 <= dataModule_io_dataOut_4_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_2 <= _GEN_4721;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_3 <= dataModule_io_dataOut_4_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_3 <= dataModule_io_dataOut_4_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_3 <= dataModule_io_dataOut_4_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_3 <= _GEN_4729;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_4 <= dataModule_io_dataOut_4_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_4 <= dataModule_io_dataOut_4_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_4 <= dataModule_io_dataOut_4_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_4 <= _GEN_4737;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_5 <= dataModule_io_dataOut_4_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_5 <= dataModule_io_dataOut_4_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_5 <= dataModule_io_dataOut_4_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_5 <= _GEN_4745;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_6 <= dataModule_io_dataOut_4_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_6 <= dataModule_io_dataOut_4_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_6 <= dataModule_io_dataOut_4_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_6 <= _GEN_4753;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_7 <= dataModule_io_dataOut_4_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_7 <= dataModule_io_dataOut_4_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__4_7 <= dataModule_io_dataOut_4_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__4_7 <= _GEN_4761;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_0 <= dataModule_io_dataOut_5_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_0 <= dataModule_io_dataOut_5_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_0 <= dataModule_io_dataOut_5_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_0 <= _GEN_4769;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_1 <= dataModule_io_dataOut_5_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_1 <= dataModule_io_dataOut_5_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_1 <= dataModule_io_dataOut_5_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_1 <= _GEN_4777;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_2 <= dataModule_io_dataOut_5_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_2 <= dataModule_io_dataOut_5_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_2 <= dataModule_io_dataOut_5_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_2 <= _GEN_4785;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_3 <= dataModule_io_dataOut_5_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_3 <= dataModule_io_dataOut_5_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_3 <= dataModule_io_dataOut_5_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_3 <= _GEN_4793;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_4 <= dataModule_io_dataOut_5_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_4 <= dataModule_io_dataOut_5_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_4 <= dataModule_io_dataOut_5_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_4 <= _GEN_4801;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_5 <= dataModule_io_dataOut_5_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_5 <= dataModule_io_dataOut_5_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_5 <= dataModule_io_dataOut_5_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_5 <= _GEN_4809;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_6 <= dataModule_io_dataOut_5_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_6 <= dataModule_io_dataOut_5_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_6 <= dataModule_io_dataOut_5_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_6 <= _GEN_4817;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_7 <= dataModule_io_dataOut_5_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_7 <= dataModule_io_dataOut_5_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__5_7 <= dataModule_io_dataOut_5_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__5_7 <= _GEN_4825;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_0 <= dataModule_io_dataOut_6_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_0 <= dataModule_io_dataOut_6_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_0 <= dataModule_io_dataOut_6_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_0 <= _GEN_4833;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_1 <= dataModule_io_dataOut_6_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_1 <= dataModule_io_dataOut_6_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_1 <= dataModule_io_dataOut_6_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_1 <= _GEN_4841;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_2 <= dataModule_io_dataOut_6_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_2 <= dataModule_io_dataOut_6_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_2 <= dataModule_io_dataOut_6_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_2 <= _GEN_4849;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_3 <= dataModule_io_dataOut_6_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_3 <= dataModule_io_dataOut_6_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_3 <= dataModule_io_dataOut_6_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_3 <= _GEN_4857;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_4 <= dataModule_io_dataOut_6_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_4 <= dataModule_io_dataOut_6_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_4 <= dataModule_io_dataOut_6_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_4 <= _GEN_4865;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_5 <= dataModule_io_dataOut_6_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_5 <= dataModule_io_dataOut_6_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_5 <= dataModule_io_dataOut_6_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_5 <= _GEN_4873;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_6 <= dataModule_io_dataOut_6_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_6 <= dataModule_io_dataOut_6_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_6 <= dataModule_io_dataOut_6_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_6 <= _GEN_4881;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_7 <= dataModule_io_dataOut_6_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_7 <= dataModule_io_dataOut_6_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__6_7 <= dataModule_io_dataOut_6_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__6_7 <= _GEN_4889;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_0 <= dataModule_io_dataOut_7_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_0 <= dataModule_io_dataOut_7_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_0 <= dataModule_io_dataOut_7_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_0 <= _GEN_4897;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_1 <= dataModule_io_dataOut_7_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_1 <= dataModule_io_dataOut_7_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_1 <= dataModule_io_dataOut_7_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_1 <= _GEN_4905;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_2 <= dataModule_io_dataOut_7_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_2 <= dataModule_io_dataOut_7_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_2 <= dataModule_io_dataOut_7_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_2 <= _GEN_4913;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_3 <= dataModule_io_dataOut_7_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_3 <= dataModule_io_dataOut_7_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_3 <= dataModule_io_dataOut_7_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_3 <= _GEN_4921;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_4 <= dataModule_io_dataOut_7_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_4 <= dataModule_io_dataOut_7_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_4 <= dataModule_io_dataOut_7_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_4 <= _GEN_4929;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_5 <= dataModule_io_dataOut_7_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_5 <= dataModule_io_dataOut_7_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_5 <= dataModule_io_dataOut_7_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_5 <= _GEN_4937;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_6 <= dataModule_io_dataOut_7_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_6 <= dataModule_io_dataOut_7_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_6 <= dataModule_io_dataOut_7_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_6 <= _GEN_4945;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_7 <= dataModule_io_dataOut_7_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_7 <= dataModule_io_dataOut_7_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__7_7 <= dataModule_io_dataOut_7_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__7_7 <= _GEN_4953;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_0 <= dataModule_io_dataOut_8_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_0 <= dataModule_io_dataOut_8_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_0 <= dataModule_io_dataOut_8_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_0 <= _GEN_4961;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_1 <= dataModule_io_dataOut_8_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_1 <= dataModule_io_dataOut_8_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_1 <= dataModule_io_dataOut_8_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_1 <= _GEN_4969;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_2 <= dataModule_io_dataOut_8_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_2 <= dataModule_io_dataOut_8_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_2 <= dataModule_io_dataOut_8_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_2 <= _GEN_4977;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_3 <= dataModule_io_dataOut_8_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_3 <= dataModule_io_dataOut_8_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_3 <= dataModule_io_dataOut_8_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_3 <= _GEN_4985;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_4 <= dataModule_io_dataOut_8_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_4 <= dataModule_io_dataOut_8_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_4 <= dataModule_io_dataOut_8_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_4 <= _GEN_4993;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_5 <= dataModule_io_dataOut_8_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_5 <= dataModule_io_dataOut_8_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_5 <= dataModule_io_dataOut_8_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_5 <= _GEN_5001;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_6 <= dataModule_io_dataOut_8_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_6 <= dataModule_io_dataOut_8_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_6 <= dataModule_io_dataOut_8_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_6 <= _GEN_5009;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_7 <= dataModule_io_dataOut_8_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_7 <= dataModule_io_dataOut_8_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__8_7 <= dataModule_io_dataOut_8_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__8_7 <= _GEN_5017;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_0 <= dataModule_io_dataOut_9_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_0 <= dataModule_io_dataOut_9_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_0 <= dataModule_io_dataOut_9_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_0 <= _GEN_5025;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_1 <= dataModule_io_dataOut_9_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_1 <= dataModule_io_dataOut_9_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_1 <= dataModule_io_dataOut_9_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_1 <= _GEN_5033;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_2 <= dataModule_io_dataOut_9_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_2 <= dataModule_io_dataOut_9_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_2 <= dataModule_io_dataOut_9_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_2 <= _GEN_5041;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_3 <= dataModule_io_dataOut_9_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_3 <= dataModule_io_dataOut_9_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_3 <= dataModule_io_dataOut_9_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_3 <= _GEN_5049;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_4 <= dataModule_io_dataOut_9_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_4 <= dataModule_io_dataOut_9_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_4 <= dataModule_io_dataOut_9_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_4 <= _GEN_5057;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_5 <= dataModule_io_dataOut_9_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_5 <= dataModule_io_dataOut_9_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_5 <= dataModule_io_dataOut_9_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_5 <= _GEN_5065;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_6 <= dataModule_io_dataOut_9_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_6 <= dataModule_io_dataOut_9_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_6 <= dataModule_io_dataOut_9_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_6 <= _GEN_5073;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_7 <= dataModule_io_dataOut_9_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_7 <= dataModule_io_dataOut_9_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__9_7 <= dataModule_io_dataOut_9_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__9_7 <= _GEN_5081;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_0 <= dataModule_io_dataOut_10_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_0 <= dataModule_io_dataOut_10_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_0 <= dataModule_io_dataOut_10_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_0 <= _GEN_5089;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_1 <= dataModule_io_dataOut_10_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_1 <= dataModule_io_dataOut_10_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_1 <= dataModule_io_dataOut_10_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_1 <= _GEN_5097;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_2 <= dataModule_io_dataOut_10_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_2 <= dataModule_io_dataOut_10_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_2 <= dataModule_io_dataOut_10_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_2 <= _GEN_5105;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_3 <= dataModule_io_dataOut_10_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_3 <= dataModule_io_dataOut_10_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_3 <= dataModule_io_dataOut_10_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_3 <= _GEN_5113;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_4 <= dataModule_io_dataOut_10_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_4 <= dataModule_io_dataOut_10_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_4 <= dataModule_io_dataOut_10_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_4 <= _GEN_5121;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_5 <= dataModule_io_dataOut_10_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_5 <= dataModule_io_dataOut_10_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_5 <= dataModule_io_dataOut_10_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_5 <= _GEN_5129;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_6 <= dataModule_io_dataOut_10_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_6 <= dataModule_io_dataOut_10_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_6 <= dataModule_io_dataOut_10_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_6 <= _GEN_5137;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_7 <= dataModule_io_dataOut_10_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_7 <= dataModule_io_dataOut_10_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__10_7 <= dataModule_io_dataOut_10_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__10_7 <= _GEN_5145;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_0 <= dataModule_io_dataOut_11_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_0 <= dataModule_io_dataOut_11_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_0 <= dataModule_io_dataOut_11_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_0 <= _GEN_5153;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_1 <= dataModule_io_dataOut_11_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_1 <= dataModule_io_dataOut_11_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_1 <= dataModule_io_dataOut_11_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_1 <= _GEN_5161;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_2 <= dataModule_io_dataOut_11_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_2 <= dataModule_io_dataOut_11_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_2 <= dataModule_io_dataOut_11_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_2 <= _GEN_5169;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_3 <= dataModule_io_dataOut_11_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_3 <= dataModule_io_dataOut_11_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_3 <= dataModule_io_dataOut_11_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_3 <= _GEN_5177;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_4 <= dataModule_io_dataOut_11_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_4 <= dataModule_io_dataOut_11_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_4 <= dataModule_io_dataOut_11_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_4 <= _GEN_5185;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_5 <= dataModule_io_dataOut_11_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_5 <= dataModule_io_dataOut_11_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_5 <= dataModule_io_dataOut_11_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_5 <= _GEN_5193;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_6 <= dataModule_io_dataOut_11_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_6 <= dataModule_io_dataOut_11_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_6 <= dataModule_io_dataOut_11_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_6 <= _GEN_5201;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_7 <= dataModule_io_dataOut_11_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_7 <= dataModule_io_dataOut_11_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__11_7 <= dataModule_io_dataOut_11_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__11_7 <= _GEN_5209;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_0 <= dataModule_io_dataOut_12_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_0 <= dataModule_io_dataOut_12_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_0 <= dataModule_io_dataOut_12_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_0 <= _GEN_5217;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_1 <= dataModule_io_dataOut_12_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_1 <= dataModule_io_dataOut_12_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_1 <= dataModule_io_dataOut_12_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_1 <= _GEN_5225;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_2 <= dataModule_io_dataOut_12_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_2 <= dataModule_io_dataOut_12_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_2 <= dataModule_io_dataOut_12_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_2 <= _GEN_5233;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_3 <= dataModule_io_dataOut_12_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_3 <= dataModule_io_dataOut_12_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_3 <= dataModule_io_dataOut_12_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_3 <= _GEN_5241;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_4 <= dataModule_io_dataOut_12_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_4 <= dataModule_io_dataOut_12_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_4 <= dataModule_io_dataOut_12_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_4 <= _GEN_5249;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_5 <= dataModule_io_dataOut_12_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_5 <= dataModule_io_dataOut_12_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_5 <= dataModule_io_dataOut_12_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_5 <= _GEN_5257;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_6 <= dataModule_io_dataOut_12_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_6 <= dataModule_io_dataOut_12_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_6 <= dataModule_io_dataOut_12_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_6 <= _GEN_5265;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_7 <= dataModule_io_dataOut_12_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_7 <= dataModule_io_dataOut_12_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__12_7 <= dataModule_io_dataOut_12_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__12_7 <= _GEN_5273;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_0 <= dataModule_io_dataOut_13_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_0 <= dataModule_io_dataOut_13_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_0 <= dataModule_io_dataOut_13_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_0 <= _GEN_5281;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_1 <= dataModule_io_dataOut_13_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_1 <= dataModule_io_dataOut_13_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_1 <= dataModule_io_dataOut_13_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_1 <= _GEN_5289;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_2 <= dataModule_io_dataOut_13_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_2 <= dataModule_io_dataOut_13_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_2 <= dataModule_io_dataOut_13_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_2 <= _GEN_5297;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_3 <= dataModule_io_dataOut_13_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_3 <= dataModule_io_dataOut_13_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_3 <= dataModule_io_dataOut_13_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_3 <= _GEN_5305;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_4 <= dataModule_io_dataOut_13_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_4 <= dataModule_io_dataOut_13_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_4 <= dataModule_io_dataOut_13_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_4 <= _GEN_5313;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_5 <= dataModule_io_dataOut_13_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_5 <= dataModule_io_dataOut_13_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_5 <= dataModule_io_dataOut_13_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_5 <= _GEN_5321;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_6 <= dataModule_io_dataOut_13_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_6 <= dataModule_io_dataOut_13_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_6 <= dataModule_io_dataOut_13_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_6 <= _GEN_5329;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_7 <= dataModule_io_dataOut_13_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_7 <= dataModule_io_dataOut_13_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__13_7 <= dataModule_io_dataOut_13_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__13_7 <= _GEN_5337;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_0 <= dataModule_io_dataOut_14_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_0 <= dataModule_io_dataOut_14_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_0 <= dataModule_io_dataOut_14_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_0 <= _GEN_5345;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_1 <= dataModule_io_dataOut_14_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_1 <= dataModule_io_dataOut_14_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_1 <= dataModule_io_dataOut_14_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_1 <= _GEN_5353;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_2 <= dataModule_io_dataOut_14_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_2 <= dataModule_io_dataOut_14_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_2 <= dataModule_io_dataOut_14_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_2 <= _GEN_5361;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_3 <= dataModule_io_dataOut_14_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_3 <= dataModule_io_dataOut_14_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_3 <= dataModule_io_dataOut_14_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_3 <= _GEN_5369;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_4 <= dataModule_io_dataOut_14_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_4 <= dataModule_io_dataOut_14_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_4 <= dataModule_io_dataOut_14_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_4 <= _GEN_5377;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_5 <= dataModule_io_dataOut_14_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_5 <= dataModule_io_dataOut_14_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_5 <= dataModule_io_dataOut_14_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_5 <= _GEN_5385;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_6 <= dataModule_io_dataOut_14_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_6 <= dataModule_io_dataOut_14_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_6 <= dataModule_io_dataOut_14_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_6 <= _GEN_5393;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_7 <= dataModule_io_dataOut_14_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_7 <= dataModule_io_dataOut_14_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__14_7 <= dataModule_io_dataOut_14_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__14_7 <= _GEN_5401;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_0 <= dataModule_io_dataOut_15_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_0 <= dataModule_io_dataOut_15_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_0 <= dataModule_io_dataOut_15_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_0 <= _GEN_5409;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_1 <= dataModule_io_dataOut_15_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_1 <= dataModule_io_dataOut_15_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_1 <= dataModule_io_dataOut_15_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_1 <= _GEN_5417;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_2 <= dataModule_io_dataOut_15_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_2 <= dataModule_io_dataOut_15_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_2 <= dataModule_io_dataOut_15_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_2 <= _GEN_5425;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_3 <= dataModule_io_dataOut_15_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_3 <= dataModule_io_dataOut_15_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_3 <= dataModule_io_dataOut_15_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_3 <= _GEN_5433;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_4 <= dataModule_io_dataOut_15_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_4 <= dataModule_io_dataOut_15_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_4 <= dataModule_io_dataOut_15_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_4 <= _GEN_5441;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_5 <= dataModule_io_dataOut_15_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_5 <= dataModule_io_dataOut_15_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_5 <= dataModule_io_dataOut_15_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_5 <= _GEN_5449;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_6 <= dataModule_io_dataOut_15_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_6 <= dataModule_io_dataOut_15_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_6 <= dataModule_io_dataOut_15_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_6 <= _GEN_5457;
      end
    end
    if (io_forward_0_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_7 <= dataModule_io_dataOut_15_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_7 <= dataModule_io_dataOut_15_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_0_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg__15_7 <= dataModule_io_dataOut_15_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg__15_7 <= _GEN_5465;
      end
    end
    valid_tag_match_reg_0_1 <= vtag_matches_1_0 & _candidateVec_T_1; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_1_1 <= vtag_matches_1_1 & _candidateVec_T_5; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_2_1 <= vtag_matches_1_2 & _candidateVec_T_9; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_3_1 <= vtag_matches_1_3 & _candidateVec_T_13; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_4_1 <= vtag_matches_1_4 & _candidateVec_T_17; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_5_1 <= vtag_matches_1_5 & _candidateVec_T_21; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_6_1 <= vtag_matches_1_6 & _candidateVec_T_25; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_7_1 <= vtag_matches_1_7 & _candidateVec_T_29; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_8_1 <= vtag_matches_1_8 & _candidateVec_T_33; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_9_1 <= vtag_matches_1_9 & _candidateVec_T_37; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_10_1 <= vtag_matches_1_10 & _candidateVec_T_41; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_11_1 <= vtag_matches_1_11 & _candidateVec_T_45; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_12_1 <= vtag_matches_1_12 & _candidateVec_T_49; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_13_1 <= vtag_matches_1_13 & _candidateVec_T_53; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_14_1 <= vtag_matches_1_14 & _candidateVec_T_57; // @[Sbuffer.scala 812:58]
    valid_tag_match_reg_15_1 <= vtag_matches_1_15 & _candidateVec_T_61; // @[Sbuffer.scala 812:58]
    inflight_tag_match_reg_0_1 <= vtag_matches_1_0 & stateVec_0_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_1_1 <= vtag_matches_1_1 & stateVec_1_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_2_1 <= vtag_matches_1_2 & stateVec_2_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_3_1 <= vtag_matches_1_3 & stateVec_3_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_4_1 <= vtag_matches_1_4 & stateVec_4_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_5_1 <= vtag_matches_1_5 & stateVec_5_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_6_1 <= vtag_matches_1_6 & stateVec_6_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_7_1 <= vtag_matches_1_7 & stateVec_7_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_8_1 <= vtag_matches_1_8 & stateVec_8_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_9_1 <= vtag_matches_1_9 & stateVec_9_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_10_1 <= vtag_matches_1_10 & stateVec_10_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_11_1 <= vtag_matches_1_11 & stateVec_11_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_12_1 <= vtag_matches_1_12 & stateVec_12_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_13_1 <= vtag_matches_1_13 & stateVec_13_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_14_1 <= vtag_matches_1_14 & stateVec_14_state_inflight; // @[Sbuffer.scala 813:61]
    inflight_tag_match_reg_15_1 <= vtag_matches_1_15 & stateVec_15_state_inflight; // @[Sbuffer.scala 813:61]
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_0 <= dataModule_io_maskOut_0_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_0 <= dataModule_io_maskOut_0_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_0 <= dataModule_io_maskOut_0_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_0 <= _GEN_5666;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_1 <= dataModule_io_maskOut_0_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_1 <= dataModule_io_maskOut_0_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_1 <= dataModule_io_maskOut_0_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_1 <= _GEN_5674;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_2 <= dataModule_io_maskOut_0_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_2 <= dataModule_io_maskOut_0_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_2 <= dataModule_io_maskOut_0_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_2 <= _GEN_5682;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_3 <= dataModule_io_maskOut_0_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_3 <= dataModule_io_maskOut_0_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_3 <= dataModule_io_maskOut_0_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_3 <= _GEN_5690;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_4 <= dataModule_io_maskOut_0_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_4 <= dataModule_io_maskOut_0_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_4 <= dataModule_io_maskOut_0_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_4 <= _GEN_5698;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_5 <= dataModule_io_maskOut_0_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_5 <= dataModule_io_maskOut_0_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_5 <= dataModule_io_maskOut_0_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_5 <= _GEN_5706;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_6 <= dataModule_io_maskOut_0_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_6 <= dataModule_io_maskOut_0_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_6 <= dataModule_io_maskOut_0_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_6 <= _GEN_5714;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_7 <= dataModule_io_maskOut_0_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_7 <= dataModule_io_maskOut_0_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_0_7 <= dataModule_io_maskOut_0_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_0_7 <= _GEN_5722;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_0 <= dataModule_io_maskOut_1_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_0 <= dataModule_io_maskOut_1_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_0 <= dataModule_io_maskOut_1_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_0 <= _GEN_5730;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_1 <= dataModule_io_maskOut_1_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_1 <= dataModule_io_maskOut_1_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_1 <= dataModule_io_maskOut_1_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_1 <= _GEN_5738;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_2 <= dataModule_io_maskOut_1_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_2 <= dataModule_io_maskOut_1_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_2 <= dataModule_io_maskOut_1_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_2 <= _GEN_5746;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_3 <= dataModule_io_maskOut_1_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_3 <= dataModule_io_maskOut_1_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_3 <= dataModule_io_maskOut_1_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_3 <= _GEN_5754;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_4 <= dataModule_io_maskOut_1_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_4 <= dataModule_io_maskOut_1_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_4 <= dataModule_io_maskOut_1_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_4 <= _GEN_5762;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_5 <= dataModule_io_maskOut_1_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_5 <= dataModule_io_maskOut_1_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_5 <= dataModule_io_maskOut_1_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_5 <= _GEN_5770;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_6 <= dataModule_io_maskOut_1_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_6 <= dataModule_io_maskOut_1_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_6 <= dataModule_io_maskOut_1_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_6 <= _GEN_5778;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_7 <= dataModule_io_maskOut_1_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_7 <= dataModule_io_maskOut_1_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_1_7 <= dataModule_io_maskOut_1_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_1_7 <= _GEN_5786;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_0 <= dataModule_io_maskOut_2_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_0 <= dataModule_io_maskOut_2_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_0 <= dataModule_io_maskOut_2_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_0 <= _GEN_5794;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_1 <= dataModule_io_maskOut_2_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_1 <= dataModule_io_maskOut_2_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_1 <= dataModule_io_maskOut_2_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_1 <= _GEN_5802;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_2 <= dataModule_io_maskOut_2_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_2 <= dataModule_io_maskOut_2_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_2 <= dataModule_io_maskOut_2_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_2 <= _GEN_5810;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_3 <= dataModule_io_maskOut_2_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_3 <= dataModule_io_maskOut_2_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_3 <= dataModule_io_maskOut_2_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_3 <= _GEN_5818;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_4 <= dataModule_io_maskOut_2_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_4 <= dataModule_io_maskOut_2_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_4 <= dataModule_io_maskOut_2_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_4 <= _GEN_5826;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_5 <= dataModule_io_maskOut_2_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_5 <= dataModule_io_maskOut_2_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_5 <= dataModule_io_maskOut_2_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_5 <= _GEN_5834;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_6 <= dataModule_io_maskOut_2_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_6 <= dataModule_io_maskOut_2_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_6 <= dataModule_io_maskOut_2_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_6 <= _GEN_5842;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_7 <= dataModule_io_maskOut_2_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_7 <= dataModule_io_maskOut_2_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_2_7 <= dataModule_io_maskOut_2_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_2_7 <= _GEN_5850;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_0 <= dataModule_io_maskOut_3_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_0 <= dataModule_io_maskOut_3_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_0 <= dataModule_io_maskOut_3_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_0 <= _GEN_5858;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_1 <= dataModule_io_maskOut_3_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_1 <= dataModule_io_maskOut_3_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_1 <= dataModule_io_maskOut_3_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_1 <= _GEN_5866;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_2 <= dataModule_io_maskOut_3_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_2 <= dataModule_io_maskOut_3_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_2 <= dataModule_io_maskOut_3_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_2 <= _GEN_5874;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_3 <= dataModule_io_maskOut_3_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_3 <= dataModule_io_maskOut_3_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_3 <= dataModule_io_maskOut_3_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_3 <= _GEN_5882;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_4 <= dataModule_io_maskOut_3_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_4 <= dataModule_io_maskOut_3_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_4 <= dataModule_io_maskOut_3_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_4 <= _GEN_5890;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_5 <= dataModule_io_maskOut_3_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_5 <= dataModule_io_maskOut_3_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_5 <= dataModule_io_maskOut_3_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_5 <= _GEN_5898;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_6 <= dataModule_io_maskOut_3_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_6 <= dataModule_io_maskOut_3_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_6 <= dataModule_io_maskOut_3_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_6 <= _GEN_5906;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_7 <= dataModule_io_maskOut_3_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_7 <= dataModule_io_maskOut_3_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_3_7 <= dataModule_io_maskOut_3_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_3_7 <= _GEN_5914;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_0 <= dataModule_io_maskOut_4_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_0 <= dataModule_io_maskOut_4_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_0 <= dataModule_io_maskOut_4_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_0 <= _GEN_5922;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_1 <= dataModule_io_maskOut_4_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_1 <= dataModule_io_maskOut_4_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_1 <= dataModule_io_maskOut_4_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_1 <= _GEN_5930;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_2 <= dataModule_io_maskOut_4_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_2 <= dataModule_io_maskOut_4_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_2 <= dataModule_io_maskOut_4_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_2 <= _GEN_5938;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_3 <= dataModule_io_maskOut_4_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_3 <= dataModule_io_maskOut_4_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_3 <= dataModule_io_maskOut_4_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_3 <= _GEN_5946;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_4 <= dataModule_io_maskOut_4_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_4 <= dataModule_io_maskOut_4_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_4 <= dataModule_io_maskOut_4_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_4 <= _GEN_5954;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_5 <= dataModule_io_maskOut_4_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_5 <= dataModule_io_maskOut_4_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_5 <= dataModule_io_maskOut_4_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_5 <= _GEN_5962;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_6 <= dataModule_io_maskOut_4_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_6 <= dataModule_io_maskOut_4_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_6 <= dataModule_io_maskOut_4_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_6 <= _GEN_5970;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_7 <= dataModule_io_maskOut_4_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_7 <= dataModule_io_maskOut_4_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_4_7 <= dataModule_io_maskOut_4_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_4_7 <= _GEN_5978;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_0 <= dataModule_io_maskOut_5_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_0 <= dataModule_io_maskOut_5_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_0 <= dataModule_io_maskOut_5_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_0 <= _GEN_5986;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_1 <= dataModule_io_maskOut_5_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_1 <= dataModule_io_maskOut_5_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_1 <= dataModule_io_maskOut_5_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_1 <= _GEN_5994;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_2 <= dataModule_io_maskOut_5_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_2 <= dataModule_io_maskOut_5_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_2 <= dataModule_io_maskOut_5_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_2 <= _GEN_6002;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_3 <= dataModule_io_maskOut_5_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_3 <= dataModule_io_maskOut_5_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_3 <= dataModule_io_maskOut_5_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_3 <= _GEN_6010;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_4 <= dataModule_io_maskOut_5_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_4 <= dataModule_io_maskOut_5_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_4 <= dataModule_io_maskOut_5_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_4 <= _GEN_6018;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_5 <= dataModule_io_maskOut_5_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_5 <= dataModule_io_maskOut_5_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_5 <= dataModule_io_maskOut_5_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_5 <= _GEN_6026;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_6 <= dataModule_io_maskOut_5_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_6 <= dataModule_io_maskOut_5_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_6 <= dataModule_io_maskOut_5_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_6 <= _GEN_6034;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_7 <= dataModule_io_maskOut_5_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_7 <= dataModule_io_maskOut_5_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_5_7 <= dataModule_io_maskOut_5_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_5_7 <= _GEN_6042;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_0 <= dataModule_io_maskOut_6_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_0 <= dataModule_io_maskOut_6_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_0 <= dataModule_io_maskOut_6_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_0 <= _GEN_6050;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_1 <= dataModule_io_maskOut_6_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_1 <= dataModule_io_maskOut_6_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_1 <= dataModule_io_maskOut_6_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_1 <= _GEN_6058;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_2 <= dataModule_io_maskOut_6_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_2 <= dataModule_io_maskOut_6_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_2 <= dataModule_io_maskOut_6_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_2 <= _GEN_6066;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_3 <= dataModule_io_maskOut_6_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_3 <= dataModule_io_maskOut_6_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_3 <= dataModule_io_maskOut_6_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_3 <= _GEN_6074;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_4 <= dataModule_io_maskOut_6_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_4 <= dataModule_io_maskOut_6_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_4 <= dataModule_io_maskOut_6_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_4 <= _GEN_6082;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_5 <= dataModule_io_maskOut_6_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_5 <= dataModule_io_maskOut_6_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_5 <= dataModule_io_maskOut_6_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_5 <= _GEN_6090;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_6 <= dataModule_io_maskOut_6_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_6 <= dataModule_io_maskOut_6_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_6 <= dataModule_io_maskOut_6_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_6 <= _GEN_6098;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_7 <= dataModule_io_maskOut_6_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_7 <= dataModule_io_maskOut_6_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_6_7 <= dataModule_io_maskOut_6_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_6_7 <= _GEN_6106;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_0 <= dataModule_io_maskOut_7_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_0 <= dataModule_io_maskOut_7_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_0 <= dataModule_io_maskOut_7_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_0 <= _GEN_6114;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_1 <= dataModule_io_maskOut_7_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_1 <= dataModule_io_maskOut_7_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_1 <= dataModule_io_maskOut_7_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_1 <= _GEN_6122;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_2 <= dataModule_io_maskOut_7_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_2 <= dataModule_io_maskOut_7_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_2 <= dataModule_io_maskOut_7_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_2 <= _GEN_6130;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_3 <= dataModule_io_maskOut_7_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_3 <= dataModule_io_maskOut_7_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_3 <= dataModule_io_maskOut_7_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_3 <= _GEN_6138;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_4 <= dataModule_io_maskOut_7_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_4 <= dataModule_io_maskOut_7_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_4 <= dataModule_io_maskOut_7_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_4 <= _GEN_6146;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_5 <= dataModule_io_maskOut_7_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_5 <= dataModule_io_maskOut_7_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_5 <= dataModule_io_maskOut_7_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_5 <= _GEN_6154;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_6 <= dataModule_io_maskOut_7_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_6 <= dataModule_io_maskOut_7_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_6 <= dataModule_io_maskOut_7_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_6 <= _GEN_6162;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_7 <= dataModule_io_maskOut_7_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_7 <= dataModule_io_maskOut_7_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_7_7 <= dataModule_io_maskOut_7_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_7_7 <= _GEN_6170;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_0 <= dataModule_io_maskOut_8_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_0 <= dataModule_io_maskOut_8_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_0 <= dataModule_io_maskOut_8_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_0 <= _GEN_6178;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_1 <= dataModule_io_maskOut_8_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_1 <= dataModule_io_maskOut_8_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_1 <= dataModule_io_maskOut_8_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_1 <= _GEN_6186;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_2 <= dataModule_io_maskOut_8_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_2 <= dataModule_io_maskOut_8_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_2 <= dataModule_io_maskOut_8_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_2 <= _GEN_6194;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_3 <= dataModule_io_maskOut_8_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_3 <= dataModule_io_maskOut_8_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_3 <= dataModule_io_maskOut_8_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_3 <= _GEN_6202;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_4 <= dataModule_io_maskOut_8_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_4 <= dataModule_io_maskOut_8_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_4 <= dataModule_io_maskOut_8_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_4 <= _GEN_6210;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_5 <= dataModule_io_maskOut_8_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_5 <= dataModule_io_maskOut_8_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_5 <= dataModule_io_maskOut_8_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_5 <= _GEN_6218;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_6 <= dataModule_io_maskOut_8_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_6 <= dataModule_io_maskOut_8_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_6 <= dataModule_io_maskOut_8_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_6 <= _GEN_6226;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_7 <= dataModule_io_maskOut_8_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_7 <= dataModule_io_maskOut_8_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_8_7 <= dataModule_io_maskOut_8_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_8_7 <= _GEN_6234;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_0 <= dataModule_io_maskOut_9_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_0 <= dataModule_io_maskOut_9_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_0 <= dataModule_io_maskOut_9_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_0 <= _GEN_6242;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_1 <= dataModule_io_maskOut_9_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_1 <= dataModule_io_maskOut_9_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_1 <= dataModule_io_maskOut_9_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_1 <= _GEN_6250;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_2 <= dataModule_io_maskOut_9_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_2 <= dataModule_io_maskOut_9_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_2 <= dataModule_io_maskOut_9_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_2 <= _GEN_6258;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_3 <= dataModule_io_maskOut_9_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_3 <= dataModule_io_maskOut_9_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_3 <= dataModule_io_maskOut_9_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_3 <= _GEN_6266;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_4 <= dataModule_io_maskOut_9_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_4 <= dataModule_io_maskOut_9_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_4 <= dataModule_io_maskOut_9_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_4 <= _GEN_6274;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_5 <= dataModule_io_maskOut_9_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_5 <= dataModule_io_maskOut_9_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_5 <= dataModule_io_maskOut_9_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_5 <= _GEN_6282;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_6 <= dataModule_io_maskOut_9_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_6 <= dataModule_io_maskOut_9_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_6 <= dataModule_io_maskOut_9_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_6 <= _GEN_6290;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_7 <= dataModule_io_maskOut_9_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_7 <= dataModule_io_maskOut_9_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_9_7 <= dataModule_io_maskOut_9_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_9_7 <= _GEN_6298;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_0 <= dataModule_io_maskOut_10_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_0 <= dataModule_io_maskOut_10_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_0 <= dataModule_io_maskOut_10_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_0 <= _GEN_6306;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_1 <= dataModule_io_maskOut_10_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_1 <= dataModule_io_maskOut_10_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_1 <= dataModule_io_maskOut_10_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_1 <= _GEN_6314;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_2 <= dataModule_io_maskOut_10_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_2 <= dataModule_io_maskOut_10_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_2 <= dataModule_io_maskOut_10_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_2 <= _GEN_6322;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_3 <= dataModule_io_maskOut_10_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_3 <= dataModule_io_maskOut_10_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_3 <= dataModule_io_maskOut_10_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_3 <= _GEN_6330;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_4 <= dataModule_io_maskOut_10_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_4 <= dataModule_io_maskOut_10_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_4 <= dataModule_io_maskOut_10_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_4 <= _GEN_6338;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_5 <= dataModule_io_maskOut_10_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_5 <= dataModule_io_maskOut_10_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_5 <= dataModule_io_maskOut_10_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_5 <= _GEN_6346;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_6 <= dataModule_io_maskOut_10_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_6 <= dataModule_io_maskOut_10_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_6 <= dataModule_io_maskOut_10_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_6 <= _GEN_6354;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_7 <= dataModule_io_maskOut_10_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_7 <= dataModule_io_maskOut_10_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_10_7 <= dataModule_io_maskOut_10_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_10_7 <= _GEN_6362;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_0 <= dataModule_io_maskOut_11_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_0 <= dataModule_io_maskOut_11_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_0 <= dataModule_io_maskOut_11_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_0 <= _GEN_6370;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_1 <= dataModule_io_maskOut_11_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_1 <= dataModule_io_maskOut_11_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_1 <= dataModule_io_maskOut_11_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_1 <= _GEN_6378;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_2 <= dataModule_io_maskOut_11_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_2 <= dataModule_io_maskOut_11_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_2 <= dataModule_io_maskOut_11_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_2 <= _GEN_6386;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_3 <= dataModule_io_maskOut_11_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_3 <= dataModule_io_maskOut_11_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_3 <= dataModule_io_maskOut_11_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_3 <= _GEN_6394;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_4 <= dataModule_io_maskOut_11_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_4 <= dataModule_io_maskOut_11_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_4 <= dataModule_io_maskOut_11_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_4 <= _GEN_6402;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_5 <= dataModule_io_maskOut_11_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_5 <= dataModule_io_maskOut_11_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_5 <= dataModule_io_maskOut_11_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_5 <= _GEN_6410;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_6 <= dataModule_io_maskOut_11_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_6 <= dataModule_io_maskOut_11_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_6 <= dataModule_io_maskOut_11_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_6 <= _GEN_6418;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_7 <= dataModule_io_maskOut_11_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_7 <= dataModule_io_maskOut_11_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_11_7 <= dataModule_io_maskOut_11_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_11_7 <= _GEN_6426;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_0 <= dataModule_io_maskOut_12_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_0 <= dataModule_io_maskOut_12_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_0 <= dataModule_io_maskOut_12_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_0 <= _GEN_6434;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_1 <= dataModule_io_maskOut_12_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_1 <= dataModule_io_maskOut_12_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_1 <= dataModule_io_maskOut_12_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_1 <= _GEN_6442;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_2 <= dataModule_io_maskOut_12_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_2 <= dataModule_io_maskOut_12_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_2 <= dataModule_io_maskOut_12_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_2 <= _GEN_6450;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_3 <= dataModule_io_maskOut_12_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_3 <= dataModule_io_maskOut_12_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_3 <= dataModule_io_maskOut_12_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_3 <= _GEN_6458;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_4 <= dataModule_io_maskOut_12_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_4 <= dataModule_io_maskOut_12_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_4 <= dataModule_io_maskOut_12_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_4 <= _GEN_6466;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_5 <= dataModule_io_maskOut_12_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_5 <= dataModule_io_maskOut_12_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_5 <= dataModule_io_maskOut_12_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_5 <= _GEN_6474;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_6 <= dataModule_io_maskOut_12_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_6 <= dataModule_io_maskOut_12_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_6 <= dataModule_io_maskOut_12_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_6 <= _GEN_6482;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_7 <= dataModule_io_maskOut_12_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_7 <= dataModule_io_maskOut_12_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_12_7 <= dataModule_io_maskOut_12_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_12_7 <= _GEN_6490;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_0 <= dataModule_io_maskOut_13_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_0 <= dataModule_io_maskOut_13_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_0 <= dataModule_io_maskOut_13_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_0 <= _GEN_6498;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_1 <= dataModule_io_maskOut_13_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_1 <= dataModule_io_maskOut_13_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_1 <= dataModule_io_maskOut_13_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_1 <= _GEN_6506;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_2 <= dataModule_io_maskOut_13_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_2 <= dataModule_io_maskOut_13_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_2 <= dataModule_io_maskOut_13_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_2 <= _GEN_6514;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_3 <= dataModule_io_maskOut_13_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_3 <= dataModule_io_maskOut_13_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_3 <= dataModule_io_maskOut_13_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_3 <= _GEN_6522;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_4 <= dataModule_io_maskOut_13_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_4 <= dataModule_io_maskOut_13_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_4 <= dataModule_io_maskOut_13_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_4 <= _GEN_6530;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_5 <= dataModule_io_maskOut_13_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_5 <= dataModule_io_maskOut_13_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_5 <= dataModule_io_maskOut_13_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_5 <= _GEN_6538;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_6 <= dataModule_io_maskOut_13_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_6 <= dataModule_io_maskOut_13_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_6 <= dataModule_io_maskOut_13_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_6 <= _GEN_6546;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_7 <= dataModule_io_maskOut_13_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_7 <= dataModule_io_maskOut_13_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_13_7 <= dataModule_io_maskOut_13_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_13_7 <= _GEN_6554;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_0 <= dataModule_io_maskOut_14_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_0 <= dataModule_io_maskOut_14_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_0 <= dataModule_io_maskOut_14_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_0 <= _GEN_6562;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_1 <= dataModule_io_maskOut_14_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_1 <= dataModule_io_maskOut_14_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_1 <= dataModule_io_maskOut_14_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_1 <= _GEN_6570;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_2 <= dataModule_io_maskOut_14_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_2 <= dataModule_io_maskOut_14_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_2 <= dataModule_io_maskOut_14_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_2 <= _GEN_6578;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_3 <= dataModule_io_maskOut_14_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_3 <= dataModule_io_maskOut_14_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_3 <= dataModule_io_maskOut_14_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_3 <= _GEN_6586;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_4 <= dataModule_io_maskOut_14_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_4 <= dataModule_io_maskOut_14_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_4 <= dataModule_io_maskOut_14_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_4 <= _GEN_6594;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_5 <= dataModule_io_maskOut_14_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_5 <= dataModule_io_maskOut_14_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_5 <= dataModule_io_maskOut_14_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_5 <= _GEN_6602;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_6 <= dataModule_io_maskOut_14_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_6 <= dataModule_io_maskOut_14_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_6 <= dataModule_io_maskOut_14_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_6 <= _GEN_6610;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_7 <= dataModule_io_maskOut_14_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_7 <= dataModule_io_maskOut_14_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_14_7 <= dataModule_io_maskOut_14_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_14_7 <= _GEN_6618;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_0 <= dataModule_io_maskOut_15_7_0; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_0 <= dataModule_io_maskOut_15_6_0; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_0 <= dataModule_io_maskOut_15_5_0; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_0 <= _GEN_6626;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_1 <= dataModule_io_maskOut_15_7_1; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_1 <= dataModule_io_maskOut_15_6_1; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_1 <= dataModule_io_maskOut_15_5_1; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_1 <= _GEN_6634;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_2 <= dataModule_io_maskOut_15_7_2; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_2 <= dataModule_io_maskOut_15_6_2; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_2 <= dataModule_io_maskOut_15_5_2; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_2 <= _GEN_6642;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_3 <= dataModule_io_maskOut_15_7_3; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_3 <= dataModule_io_maskOut_15_6_3; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_3 <= dataModule_io_maskOut_15_5_3; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_3 <= _GEN_6650;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_4 <= dataModule_io_maskOut_15_7_4; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_4 <= dataModule_io_maskOut_15_6_4; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_4 <= dataModule_io_maskOut_15_5_4; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_4 <= _GEN_6658;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_5 <= dataModule_io_maskOut_15_7_5; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_5 <= dataModule_io_maskOut_15_6_5; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_5 <= dataModule_io_maskOut_15_5_5; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_5 <= _GEN_6666;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_6 <= dataModule_io_maskOut_15_7_6; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_6 <= dataModule_io_maskOut_15_6_6; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_6 <= dataModule_io_maskOut_15_5_6; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_6 <= _GEN_6674;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_7 <= dataModule_io_maskOut_15_7_7; // @[Sbuffer.scala 820:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_7 <= dataModule_io_maskOut_15_6_7; // @[Sbuffer.scala 820:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 820:14]
        forward_mask_candidate_reg_1_15_7 <= dataModule_io_maskOut_15_5_7; // @[Sbuffer.scala 820:14]
      end else begin
        forward_mask_candidate_reg_1_15_7 <= _GEN_6682;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_0 <= dataModule_io_dataOut_0_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_0 <= dataModule_io_dataOut_0_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_0 <= dataModule_io_dataOut_0_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_0 <= _GEN_6818;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_1 <= dataModule_io_dataOut_0_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_1 <= dataModule_io_dataOut_0_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_1 <= dataModule_io_dataOut_0_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_1 <= _GEN_6826;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_2 <= dataModule_io_dataOut_0_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_2 <= dataModule_io_dataOut_0_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_2 <= dataModule_io_dataOut_0_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_2 <= _GEN_6834;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_3 <= dataModule_io_dataOut_0_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_3 <= dataModule_io_dataOut_0_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_3 <= dataModule_io_dataOut_0_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_3 <= _GEN_6842;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_4 <= dataModule_io_dataOut_0_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_4 <= dataModule_io_dataOut_0_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_4 <= dataModule_io_dataOut_0_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_4 <= _GEN_6850;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_5 <= dataModule_io_dataOut_0_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_5 <= dataModule_io_dataOut_0_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_5 <= dataModule_io_dataOut_0_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_5 <= _GEN_6858;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_6 <= dataModule_io_dataOut_0_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_6 <= dataModule_io_dataOut_0_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_6 <= dataModule_io_dataOut_0_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_6 <= _GEN_6866;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_7 <= dataModule_io_dataOut_0_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_7 <= dataModule_io_dataOut_0_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_0_7 <= dataModule_io_dataOut_0_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_0_7 <= _GEN_6874;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_0 <= dataModule_io_dataOut_1_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_0 <= dataModule_io_dataOut_1_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_0 <= dataModule_io_dataOut_1_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_0 <= _GEN_6882;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_1 <= dataModule_io_dataOut_1_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_1 <= dataModule_io_dataOut_1_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_1 <= dataModule_io_dataOut_1_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_1 <= _GEN_6890;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_2 <= dataModule_io_dataOut_1_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_2 <= dataModule_io_dataOut_1_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_2 <= dataModule_io_dataOut_1_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_2 <= _GEN_6898;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_3 <= dataModule_io_dataOut_1_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_3 <= dataModule_io_dataOut_1_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_3 <= dataModule_io_dataOut_1_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_3 <= _GEN_6906;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_4 <= dataModule_io_dataOut_1_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_4 <= dataModule_io_dataOut_1_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_4 <= dataModule_io_dataOut_1_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_4 <= _GEN_6914;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_5 <= dataModule_io_dataOut_1_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_5 <= dataModule_io_dataOut_1_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_5 <= dataModule_io_dataOut_1_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_5 <= _GEN_6922;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_6 <= dataModule_io_dataOut_1_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_6 <= dataModule_io_dataOut_1_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_6 <= dataModule_io_dataOut_1_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_6 <= _GEN_6930;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_7 <= dataModule_io_dataOut_1_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_7 <= dataModule_io_dataOut_1_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_1_7 <= dataModule_io_dataOut_1_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_1_7 <= _GEN_6938;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_0 <= dataModule_io_dataOut_2_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_0 <= dataModule_io_dataOut_2_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_0 <= dataModule_io_dataOut_2_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_0 <= _GEN_6946;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_1 <= dataModule_io_dataOut_2_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_1 <= dataModule_io_dataOut_2_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_1 <= dataModule_io_dataOut_2_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_1 <= _GEN_6954;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_2 <= dataModule_io_dataOut_2_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_2 <= dataModule_io_dataOut_2_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_2 <= dataModule_io_dataOut_2_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_2 <= _GEN_6962;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_3 <= dataModule_io_dataOut_2_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_3 <= dataModule_io_dataOut_2_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_3 <= dataModule_io_dataOut_2_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_3 <= _GEN_6970;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_4 <= dataModule_io_dataOut_2_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_4 <= dataModule_io_dataOut_2_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_4 <= dataModule_io_dataOut_2_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_4 <= _GEN_6978;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_5 <= dataModule_io_dataOut_2_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_5 <= dataModule_io_dataOut_2_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_5 <= dataModule_io_dataOut_2_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_5 <= _GEN_6986;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_6 <= dataModule_io_dataOut_2_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_6 <= dataModule_io_dataOut_2_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_6 <= dataModule_io_dataOut_2_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_6 <= _GEN_6994;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_7 <= dataModule_io_dataOut_2_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_7 <= dataModule_io_dataOut_2_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_2_7 <= dataModule_io_dataOut_2_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_2_7 <= _GEN_7002;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_0 <= dataModule_io_dataOut_3_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_0 <= dataModule_io_dataOut_3_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_0 <= dataModule_io_dataOut_3_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_0 <= _GEN_7010;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_1 <= dataModule_io_dataOut_3_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_1 <= dataModule_io_dataOut_3_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_1 <= dataModule_io_dataOut_3_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_1 <= _GEN_7018;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_2 <= dataModule_io_dataOut_3_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_2 <= dataModule_io_dataOut_3_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_2 <= dataModule_io_dataOut_3_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_2 <= _GEN_7026;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_3 <= dataModule_io_dataOut_3_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_3 <= dataModule_io_dataOut_3_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_3 <= dataModule_io_dataOut_3_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_3 <= _GEN_7034;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_4 <= dataModule_io_dataOut_3_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_4 <= dataModule_io_dataOut_3_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_4 <= dataModule_io_dataOut_3_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_4 <= _GEN_7042;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_5 <= dataModule_io_dataOut_3_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_5 <= dataModule_io_dataOut_3_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_5 <= dataModule_io_dataOut_3_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_5 <= _GEN_7050;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_6 <= dataModule_io_dataOut_3_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_6 <= dataModule_io_dataOut_3_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_6 <= dataModule_io_dataOut_3_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_6 <= _GEN_7058;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_7 <= dataModule_io_dataOut_3_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_7 <= dataModule_io_dataOut_3_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_3_7 <= dataModule_io_dataOut_3_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_3_7 <= _GEN_7066;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_0 <= dataModule_io_dataOut_4_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_0 <= dataModule_io_dataOut_4_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_0 <= dataModule_io_dataOut_4_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_0 <= _GEN_7074;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_1 <= dataModule_io_dataOut_4_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_1 <= dataModule_io_dataOut_4_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_1 <= dataModule_io_dataOut_4_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_1 <= _GEN_7082;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_2 <= dataModule_io_dataOut_4_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_2 <= dataModule_io_dataOut_4_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_2 <= dataModule_io_dataOut_4_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_2 <= _GEN_7090;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_3 <= dataModule_io_dataOut_4_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_3 <= dataModule_io_dataOut_4_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_3 <= dataModule_io_dataOut_4_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_3 <= _GEN_7098;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_4 <= dataModule_io_dataOut_4_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_4 <= dataModule_io_dataOut_4_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_4 <= dataModule_io_dataOut_4_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_4 <= _GEN_7106;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_5 <= dataModule_io_dataOut_4_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_5 <= dataModule_io_dataOut_4_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_5 <= dataModule_io_dataOut_4_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_5 <= _GEN_7114;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_6 <= dataModule_io_dataOut_4_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_6 <= dataModule_io_dataOut_4_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_6 <= dataModule_io_dataOut_4_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_6 <= _GEN_7122;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_7 <= dataModule_io_dataOut_4_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_7 <= dataModule_io_dataOut_4_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_4_7 <= dataModule_io_dataOut_4_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_4_7 <= _GEN_7130;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_0 <= dataModule_io_dataOut_5_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_0 <= dataModule_io_dataOut_5_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_0 <= dataModule_io_dataOut_5_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_0 <= _GEN_7138;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_1 <= dataModule_io_dataOut_5_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_1 <= dataModule_io_dataOut_5_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_1 <= dataModule_io_dataOut_5_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_1 <= _GEN_7146;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_2 <= dataModule_io_dataOut_5_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_2 <= dataModule_io_dataOut_5_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_2 <= dataModule_io_dataOut_5_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_2 <= _GEN_7154;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_3 <= dataModule_io_dataOut_5_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_3 <= dataModule_io_dataOut_5_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_3 <= dataModule_io_dataOut_5_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_3 <= _GEN_7162;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_4 <= dataModule_io_dataOut_5_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_4 <= dataModule_io_dataOut_5_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_4 <= dataModule_io_dataOut_5_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_4 <= _GEN_7170;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_5 <= dataModule_io_dataOut_5_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_5 <= dataModule_io_dataOut_5_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_5 <= dataModule_io_dataOut_5_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_5 <= _GEN_7178;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_6 <= dataModule_io_dataOut_5_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_6 <= dataModule_io_dataOut_5_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_6 <= dataModule_io_dataOut_5_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_6 <= _GEN_7186;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_7 <= dataModule_io_dataOut_5_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_7 <= dataModule_io_dataOut_5_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_5_7 <= dataModule_io_dataOut_5_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_5_7 <= _GEN_7194;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_0 <= dataModule_io_dataOut_6_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_0 <= dataModule_io_dataOut_6_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_0 <= dataModule_io_dataOut_6_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_0 <= _GEN_7202;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_1 <= dataModule_io_dataOut_6_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_1 <= dataModule_io_dataOut_6_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_1 <= dataModule_io_dataOut_6_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_1 <= _GEN_7210;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_2 <= dataModule_io_dataOut_6_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_2 <= dataModule_io_dataOut_6_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_2 <= dataModule_io_dataOut_6_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_2 <= _GEN_7218;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_3 <= dataModule_io_dataOut_6_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_3 <= dataModule_io_dataOut_6_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_3 <= dataModule_io_dataOut_6_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_3 <= _GEN_7226;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_4 <= dataModule_io_dataOut_6_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_4 <= dataModule_io_dataOut_6_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_4 <= dataModule_io_dataOut_6_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_4 <= _GEN_7234;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_5 <= dataModule_io_dataOut_6_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_5 <= dataModule_io_dataOut_6_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_5 <= dataModule_io_dataOut_6_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_5 <= _GEN_7242;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_6 <= dataModule_io_dataOut_6_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_6 <= dataModule_io_dataOut_6_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_6 <= dataModule_io_dataOut_6_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_6 <= _GEN_7250;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_7 <= dataModule_io_dataOut_6_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_7 <= dataModule_io_dataOut_6_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_6_7 <= dataModule_io_dataOut_6_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_6_7 <= _GEN_7258;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_0 <= dataModule_io_dataOut_7_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_0 <= dataModule_io_dataOut_7_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_0 <= dataModule_io_dataOut_7_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_0 <= _GEN_7266;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_1 <= dataModule_io_dataOut_7_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_1 <= dataModule_io_dataOut_7_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_1 <= dataModule_io_dataOut_7_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_1 <= _GEN_7274;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_2 <= dataModule_io_dataOut_7_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_2 <= dataModule_io_dataOut_7_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_2 <= dataModule_io_dataOut_7_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_2 <= _GEN_7282;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_3 <= dataModule_io_dataOut_7_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_3 <= dataModule_io_dataOut_7_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_3 <= dataModule_io_dataOut_7_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_3 <= _GEN_7290;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_4 <= dataModule_io_dataOut_7_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_4 <= dataModule_io_dataOut_7_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_4 <= dataModule_io_dataOut_7_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_4 <= _GEN_7298;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_5 <= dataModule_io_dataOut_7_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_5 <= dataModule_io_dataOut_7_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_5 <= dataModule_io_dataOut_7_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_5 <= _GEN_7306;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_6 <= dataModule_io_dataOut_7_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_6 <= dataModule_io_dataOut_7_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_6 <= dataModule_io_dataOut_7_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_6 <= _GEN_7314;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_7 <= dataModule_io_dataOut_7_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_7 <= dataModule_io_dataOut_7_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_7_7 <= dataModule_io_dataOut_7_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_7_7 <= _GEN_7322;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_0 <= dataModule_io_dataOut_8_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_0 <= dataModule_io_dataOut_8_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_0 <= dataModule_io_dataOut_8_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_0 <= _GEN_7330;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_1 <= dataModule_io_dataOut_8_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_1 <= dataModule_io_dataOut_8_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_1 <= dataModule_io_dataOut_8_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_1 <= _GEN_7338;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_2 <= dataModule_io_dataOut_8_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_2 <= dataModule_io_dataOut_8_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_2 <= dataModule_io_dataOut_8_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_2 <= _GEN_7346;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_3 <= dataModule_io_dataOut_8_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_3 <= dataModule_io_dataOut_8_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_3 <= dataModule_io_dataOut_8_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_3 <= _GEN_7354;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_4 <= dataModule_io_dataOut_8_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_4 <= dataModule_io_dataOut_8_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_4 <= dataModule_io_dataOut_8_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_4 <= _GEN_7362;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_5 <= dataModule_io_dataOut_8_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_5 <= dataModule_io_dataOut_8_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_5 <= dataModule_io_dataOut_8_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_5 <= _GEN_7370;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_6 <= dataModule_io_dataOut_8_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_6 <= dataModule_io_dataOut_8_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_6 <= dataModule_io_dataOut_8_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_6 <= _GEN_7378;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_7 <= dataModule_io_dataOut_8_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_7 <= dataModule_io_dataOut_8_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_8_7 <= dataModule_io_dataOut_8_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_8_7 <= _GEN_7386;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_0 <= dataModule_io_dataOut_9_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_0 <= dataModule_io_dataOut_9_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_0 <= dataModule_io_dataOut_9_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_0 <= _GEN_7394;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_1 <= dataModule_io_dataOut_9_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_1 <= dataModule_io_dataOut_9_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_1 <= dataModule_io_dataOut_9_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_1 <= _GEN_7402;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_2 <= dataModule_io_dataOut_9_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_2 <= dataModule_io_dataOut_9_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_2 <= dataModule_io_dataOut_9_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_2 <= _GEN_7410;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_3 <= dataModule_io_dataOut_9_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_3 <= dataModule_io_dataOut_9_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_3 <= dataModule_io_dataOut_9_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_3 <= _GEN_7418;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_4 <= dataModule_io_dataOut_9_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_4 <= dataModule_io_dataOut_9_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_4 <= dataModule_io_dataOut_9_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_4 <= _GEN_7426;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_5 <= dataModule_io_dataOut_9_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_5 <= dataModule_io_dataOut_9_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_5 <= dataModule_io_dataOut_9_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_5 <= _GEN_7434;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_6 <= dataModule_io_dataOut_9_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_6 <= dataModule_io_dataOut_9_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_6 <= dataModule_io_dataOut_9_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_6 <= _GEN_7442;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_7 <= dataModule_io_dataOut_9_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_7 <= dataModule_io_dataOut_9_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_9_7 <= dataModule_io_dataOut_9_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_9_7 <= _GEN_7450;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_0 <= dataModule_io_dataOut_10_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_0 <= dataModule_io_dataOut_10_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_0 <= dataModule_io_dataOut_10_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_0 <= _GEN_7458;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_1 <= dataModule_io_dataOut_10_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_1 <= dataModule_io_dataOut_10_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_1 <= dataModule_io_dataOut_10_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_1 <= _GEN_7466;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_2 <= dataModule_io_dataOut_10_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_2 <= dataModule_io_dataOut_10_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_2 <= dataModule_io_dataOut_10_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_2 <= _GEN_7474;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_3 <= dataModule_io_dataOut_10_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_3 <= dataModule_io_dataOut_10_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_3 <= dataModule_io_dataOut_10_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_3 <= _GEN_7482;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_4 <= dataModule_io_dataOut_10_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_4 <= dataModule_io_dataOut_10_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_4 <= dataModule_io_dataOut_10_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_4 <= _GEN_7490;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_5 <= dataModule_io_dataOut_10_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_5 <= dataModule_io_dataOut_10_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_5 <= dataModule_io_dataOut_10_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_5 <= _GEN_7498;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_6 <= dataModule_io_dataOut_10_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_6 <= dataModule_io_dataOut_10_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_6 <= dataModule_io_dataOut_10_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_6 <= _GEN_7506;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_7 <= dataModule_io_dataOut_10_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_7 <= dataModule_io_dataOut_10_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_10_7 <= dataModule_io_dataOut_10_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_10_7 <= _GEN_7514;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_0 <= dataModule_io_dataOut_11_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_0 <= dataModule_io_dataOut_11_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_0 <= dataModule_io_dataOut_11_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_0 <= _GEN_7522;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_1 <= dataModule_io_dataOut_11_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_1 <= dataModule_io_dataOut_11_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_1 <= dataModule_io_dataOut_11_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_1 <= _GEN_7530;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_2 <= dataModule_io_dataOut_11_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_2 <= dataModule_io_dataOut_11_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_2 <= dataModule_io_dataOut_11_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_2 <= _GEN_7538;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_3 <= dataModule_io_dataOut_11_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_3 <= dataModule_io_dataOut_11_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_3 <= dataModule_io_dataOut_11_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_3 <= _GEN_7546;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_4 <= dataModule_io_dataOut_11_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_4 <= dataModule_io_dataOut_11_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_4 <= dataModule_io_dataOut_11_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_4 <= _GEN_7554;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_5 <= dataModule_io_dataOut_11_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_5 <= dataModule_io_dataOut_11_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_5 <= dataModule_io_dataOut_11_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_5 <= _GEN_7562;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_6 <= dataModule_io_dataOut_11_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_6 <= dataModule_io_dataOut_11_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_6 <= dataModule_io_dataOut_11_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_6 <= _GEN_7570;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_7 <= dataModule_io_dataOut_11_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_7 <= dataModule_io_dataOut_11_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_11_7 <= dataModule_io_dataOut_11_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_11_7 <= _GEN_7578;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_0 <= dataModule_io_dataOut_12_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_0 <= dataModule_io_dataOut_12_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_0 <= dataModule_io_dataOut_12_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_0 <= _GEN_7586;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_1 <= dataModule_io_dataOut_12_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_1 <= dataModule_io_dataOut_12_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_1 <= dataModule_io_dataOut_12_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_1 <= _GEN_7594;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_2 <= dataModule_io_dataOut_12_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_2 <= dataModule_io_dataOut_12_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_2 <= dataModule_io_dataOut_12_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_2 <= _GEN_7602;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_3 <= dataModule_io_dataOut_12_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_3 <= dataModule_io_dataOut_12_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_3 <= dataModule_io_dataOut_12_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_3 <= _GEN_7610;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_4 <= dataModule_io_dataOut_12_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_4 <= dataModule_io_dataOut_12_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_4 <= dataModule_io_dataOut_12_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_4 <= _GEN_7618;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_5 <= dataModule_io_dataOut_12_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_5 <= dataModule_io_dataOut_12_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_5 <= dataModule_io_dataOut_12_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_5 <= _GEN_7626;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_6 <= dataModule_io_dataOut_12_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_6 <= dataModule_io_dataOut_12_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_6 <= dataModule_io_dataOut_12_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_6 <= _GEN_7634;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_7 <= dataModule_io_dataOut_12_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_7 <= dataModule_io_dataOut_12_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_12_7 <= dataModule_io_dataOut_12_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_12_7 <= _GEN_7642;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_0 <= dataModule_io_dataOut_13_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_0 <= dataModule_io_dataOut_13_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_0 <= dataModule_io_dataOut_13_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_0 <= _GEN_7650;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_1 <= dataModule_io_dataOut_13_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_1 <= dataModule_io_dataOut_13_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_1 <= dataModule_io_dataOut_13_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_1 <= _GEN_7658;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_2 <= dataModule_io_dataOut_13_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_2 <= dataModule_io_dataOut_13_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_2 <= dataModule_io_dataOut_13_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_2 <= _GEN_7666;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_3 <= dataModule_io_dataOut_13_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_3 <= dataModule_io_dataOut_13_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_3 <= dataModule_io_dataOut_13_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_3 <= _GEN_7674;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_4 <= dataModule_io_dataOut_13_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_4 <= dataModule_io_dataOut_13_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_4 <= dataModule_io_dataOut_13_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_4 <= _GEN_7682;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_5 <= dataModule_io_dataOut_13_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_5 <= dataModule_io_dataOut_13_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_5 <= dataModule_io_dataOut_13_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_5 <= _GEN_7690;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_6 <= dataModule_io_dataOut_13_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_6 <= dataModule_io_dataOut_13_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_6 <= dataModule_io_dataOut_13_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_6 <= _GEN_7698;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_7 <= dataModule_io_dataOut_13_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_7 <= dataModule_io_dataOut_13_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_13_7 <= dataModule_io_dataOut_13_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_13_7 <= _GEN_7706;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_0 <= dataModule_io_dataOut_14_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_0 <= dataModule_io_dataOut_14_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_0 <= dataModule_io_dataOut_14_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_0 <= _GEN_7714;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_1 <= dataModule_io_dataOut_14_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_1 <= dataModule_io_dataOut_14_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_1 <= dataModule_io_dataOut_14_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_1 <= _GEN_7722;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_2 <= dataModule_io_dataOut_14_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_2 <= dataModule_io_dataOut_14_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_2 <= dataModule_io_dataOut_14_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_2 <= _GEN_7730;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_3 <= dataModule_io_dataOut_14_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_3 <= dataModule_io_dataOut_14_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_3 <= dataModule_io_dataOut_14_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_3 <= _GEN_7738;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_4 <= dataModule_io_dataOut_14_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_4 <= dataModule_io_dataOut_14_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_4 <= dataModule_io_dataOut_14_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_4 <= _GEN_7746;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_5 <= dataModule_io_dataOut_14_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_5 <= dataModule_io_dataOut_14_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_5 <= dataModule_io_dataOut_14_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_5 <= _GEN_7754;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_6 <= dataModule_io_dataOut_14_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_6 <= dataModule_io_dataOut_14_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_6 <= dataModule_io_dataOut_14_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_6 <= _GEN_7762;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_7 <= dataModule_io_dataOut_14_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_7 <= dataModule_io_dataOut_14_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_14_7 <= dataModule_io_dataOut_14_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_14_7 <= _GEN_7770;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_0 <= dataModule_io_dataOut_15_7_0; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_0 <= dataModule_io_dataOut_15_6_0; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_0 <= dataModule_io_dataOut_15_5_0; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_0 <= _GEN_7778;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_1 <= dataModule_io_dataOut_15_7_1; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_1 <= dataModule_io_dataOut_15_6_1; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_1 <= dataModule_io_dataOut_15_5_1; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_1 <= _GEN_7786;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_2 <= dataModule_io_dataOut_15_7_2; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_2 <= dataModule_io_dataOut_15_6_2; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_2 <= dataModule_io_dataOut_15_5_2; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_2 <= _GEN_7794;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_3 <= dataModule_io_dataOut_15_7_3; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_3 <= dataModule_io_dataOut_15_6_3; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_3 <= dataModule_io_dataOut_15_5_3; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_3 <= _GEN_7802;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_4 <= dataModule_io_dataOut_15_7_4; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_4 <= dataModule_io_dataOut_15_6_4; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_4 <= dataModule_io_dataOut_15_5_4; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_4 <= _GEN_7810;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_5 <= dataModule_io_dataOut_15_7_5; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_5 <= dataModule_io_dataOut_15_6_5; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_5 <= dataModule_io_dataOut_15_5_5; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_5 <= _GEN_7818;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_6 <= dataModule_io_dataOut_15_7_6; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_6 <= dataModule_io_dataOut_15_6_6; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_6 <= dataModule_io_dataOut_15_5_6; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_6 <= _GEN_7826;
      end
    end
    if (io_forward_1_valid) begin // @[Reg.scala 20:18]
      if (3'h7 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_7 <= dataModule_io_dataOut_15_7_7; // @[Sbuffer.scala 824:14]
      end else if (3'h6 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_7 <= dataModule_io_dataOut_15_6_7; // @[Sbuffer.scala 824:14]
      end else if (3'h5 == io_forward_1_paddr[5:3]) begin // @[Sbuffer.scala 824:14]
        forward_data_candidate_reg_1_15_7 <= dataModule_io_dataOut_15_5_7; // @[Sbuffer.scala 824:14]
      end else begin
        forward_data_candidate_reg_1_15_7 <= _GEN_7834;
      end
    end
    perf_valid_entry_count <= _perf_valid_entry_count_T_61 + _perf_valid_entry_count_T_75; // @[Bitwise.scala 51:90]
    io_perf_0_value_REG <= _T_1099[0] + _T_1099[1]; // @[Bitwise.scala 51:90]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_1_value_REG <= _T_1106[0] + _T_1106[1]; // @[Bitwise.scala 51:90]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_2_value_REG <= _T_1115[0] + _T_1115[1]; // @[Bitwise.scala 51:90]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_3_value_REG <= _T_1126[0] + _T_1126[1]; // @[Bitwise.scala 51:90]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_4_value_REG <= io_dcache_req_valid; // @[PerfCounterUtils.scala 172:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_5_value_REG <= io_dcache_req_ready & io_dcache_req_valid; // @[Decoupled.scala 51:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_6_value_REG <= sbuffer_state == 2'h0; // @[Sbuffer.scala 902:42]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_7_value_REG <= sbuffer_state == 2'h3; // @[Sbuffer.scala 903:42]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_8_value_REG <= sbuffer_state == 2'h1; // @[Sbuffer.scala 904:42]
    io_perf_8_value_REG_1 <= io_perf_8_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_9_value_REG <= io_dcache_main_pipe_hit_resp_valid; // @[PerfCounterUtils.scala 172:35]
    io_perf_9_value_REG_1 <= io_perf_9_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_10_value_REG <= io_dcache_refill_hit_resp_valid; // @[PerfCounterUtils.scala 172:35]
    io_perf_10_value_REG_1 <= io_perf_10_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_11_value_REG <= io_dcache_replay_resp_valid; // @[PerfCounterUtils.scala 172:35]
    io_perf_11_value_REG_1 <= io_perf_11_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_12_value_REG <= cohTimeOutMask_0 | f_tail_13; // @[PriorityMuxDefault.scala 46:46]
    io_perf_12_value_REG_1 <= io_perf_12_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_13_value_REG <= perf_valid_entry_count < _T_1135; // @[Sbuffer.scala 909:52]
    io_perf_13_value_REG_1 <= io_perf_13_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_14_value_REG <= perf_valid_entry_count > _T_1135 & perf_valid_entry_count <= _T_1139; // @[Sbuffer.scala 910:79]
    io_perf_14_value_REG_1 <= io_perf_14_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_15_value_REG <= perf_valid_entry_count > _T_1139 & _GEN_3180 <= _T_1145; // @[Sbuffer.scala 911:79]
    io_perf_15_value_REG_1 <= io_perf_15_value_REG; // @[PerfCounterUtils.scala 172:27]
    io_perf_16_value_REG <= _GEN_3180 > _T_1145; // @[Sbuffer.scala 912:52]
    io_perf_16_value_REG_1 <= io_perf_16_value_REG; // @[PerfCounterUtils.scala 172:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_0_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h0 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_0_state_valid <= 1'h0;
      end else begin
        stateVec_0_state_valid <= _GEN_3020;
      end
    end else begin
      stateVec_0_state_valid <= _GEN_3020;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_0_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h0 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_0_state_inflight <= 1'h0;
      end else begin
        stateVec_0_state_inflight <= _GEN_3004;
      end
    end else begin
      stateVec_0_state_inflight <= _GEN_3004;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_0_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_0_w_timeout <= _GEN_3164; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h0 == sbuffer_out_s0_evictionIdx) begin
        stateVec_0_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_0_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_829) begin // @[Sbuffer.scala 745:8]
      stateVec_0_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_718) begin // @[Sbuffer.scala 511:20]
      stateVec_0_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_0_w_sameblock_inflight <= _GEN_279;
      end else begin
        stateVec_0_w_sameblock_inflight <= _GEN_408;
      end
    end else begin
      stateVec_0_w_sameblock_inflight <= _GEN_279;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_1_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h1 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_1_state_valid <= 1'h0;
      end else begin
        stateVec_1_state_valid <= _GEN_3021;
      end
    end else begin
      stateVec_1_state_valid <= _GEN_3021;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_1_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h1 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_1_state_inflight <= 1'h0;
      end else begin
        stateVec_1_state_inflight <= _GEN_3005;
      end
    end else begin
      stateVec_1_state_inflight <= _GEN_3005;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_1_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_1_w_timeout <= _GEN_3165; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h1 == sbuffer_out_s0_evictionIdx) begin
        stateVec_1_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_1_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_835) begin // @[Sbuffer.scala 745:8]
      stateVec_1_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_724) begin // @[Sbuffer.scala 511:20]
      stateVec_1_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_1_w_sameblock_inflight <= _GEN_284;
      end else begin
        stateVec_1_w_sameblock_inflight <= _GEN_415;
      end
    end else begin
      stateVec_1_w_sameblock_inflight <= _GEN_284;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_2_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h2 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_2_state_valid <= 1'h0;
      end else begin
        stateVec_2_state_valid <= _GEN_3022;
      end
    end else begin
      stateVec_2_state_valid <= _GEN_3022;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_2_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h2 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_2_state_inflight <= 1'h0;
      end else begin
        stateVec_2_state_inflight <= _GEN_3006;
      end
    end else begin
      stateVec_2_state_inflight <= _GEN_3006;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_2_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_2_w_timeout <= _GEN_3166; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h2 == sbuffer_out_s0_evictionIdx) begin
        stateVec_2_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_2_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_841) begin // @[Sbuffer.scala 745:8]
      stateVec_2_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_730) begin // @[Sbuffer.scala 511:20]
      stateVec_2_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_2_w_sameblock_inflight <= _GEN_289;
      end else begin
        stateVec_2_w_sameblock_inflight <= _GEN_422;
      end
    end else begin
      stateVec_2_w_sameblock_inflight <= _GEN_289;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_3_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h3 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_3_state_valid <= 1'h0;
      end else begin
        stateVec_3_state_valid <= _GEN_3023;
      end
    end else begin
      stateVec_3_state_valid <= _GEN_3023;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_3_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h3 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_3_state_inflight <= 1'h0;
      end else begin
        stateVec_3_state_inflight <= _GEN_3007;
      end
    end else begin
      stateVec_3_state_inflight <= _GEN_3007;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_3_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_3_w_timeout <= _GEN_3167; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h3 == sbuffer_out_s0_evictionIdx) begin
        stateVec_3_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_3_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_847) begin // @[Sbuffer.scala 745:8]
      stateVec_3_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_736) begin // @[Sbuffer.scala 511:20]
      stateVec_3_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_3_w_sameblock_inflight <= _GEN_294;
      end else begin
        stateVec_3_w_sameblock_inflight <= _GEN_429;
      end
    end else begin
      stateVec_3_w_sameblock_inflight <= _GEN_294;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_4_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h4 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_4_state_valid <= 1'h0;
      end else begin
        stateVec_4_state_valid <= _GEN_3024;
      end
    end else begin
      stateVec_4_state_valid <= _GEN_3024;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_4_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h4 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_4_state_inflight <= 1'h0;
      end else begin
        stateVec_4_state_inflight <= _GEN_3008;
      end
    end else begin
      stateVec_4_state_inflight <= _GEN_3008;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_4_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_4_w_timeout <= _GEN_3168; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h4 == sbuffer_out_s0_evictionIdx) begin
        stateVec_4_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_4_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_853) begin // @[Sbuffer.scala 745:8]
      stateVec_4_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_742) begin // @[Sbuffer.scala 511:20]
      stateVec_4_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_4_w_sameblock_inflight <= _GEN_299;
      end else begin
        stateVec_4_w_sameblock_inflight <= _GEN_436;
      end
    end else begin
      stateVec_4_w_sameblock_inflight <= _GEN_299;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_5_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h5 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_5_state_valid <= 1'h0;
      end else begin
        stateVec_5_state_valid <= _GEN_3025;
      end
    end else begin
      stateVec_5_state_valid <= _GEN_3025;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_5_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h5 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_5_state_inflight <= 1'h0;
      end else begin
        stateVec_5_state_inflight <= _GEN_3009;
      end
    end else begin
      stateVec_5_state_inflight <= _GEN_3009;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_5_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_5_w_timeout <= _GEN_3169; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h5 == sbuffer_out_s0_evictionIdx) begin
        stateVec_5_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_5_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_859) begin // @[Sbuffer.scala 745:8]
      stateVec_5_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_748) begin // @[Sbuffer.scala 511:20]
      stateVec_5_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_5_w_sameblock_inflight <= _GEN_304;
      end else begin
        stateVec_5_w_sameblock_inflight <= _GEN_443;
      end
    end else begin
      stateVec_5_w_sameblock_inflight <= _GEN_304;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_6_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h6 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_6_state_valid <= 1'h0;
      end else begin
        stateVec_6_state_valid <= _GEN_3026;
      end
    end else begin
      stateVec_6_state_valid <= _GEN_3026;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_6_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h6 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_6_state_inflight <= 1'h0;
      end else begin
        stateVec_6_state_inflight <= _GEN_3010;
      end
    end else begin
      stateVec_6_state_inflight <= _GEN_3010;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_6_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_6_w_timeout <= _GEN_3170; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h6 == sbuffer_out_s0_evictionIdx) begin
        stateVec_6_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_6_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_865) begin // @[Sbuffer.scala 745:8]
      stateVec_6_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_754) begin // @[Sbuffer.scala 511:20]
      stateVec_6_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_6_w_sameblock_inflight <= _GEN_309;
      end else begin
        stateVec_6_w_sameblock_inflight <= _GEN_450;
      end
    end else begin
      stateVec_6_w_sameblock_inflight <= _GEN_309;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_7_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h7 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_7_state_valid <= 1'h0;
      end else begin
        stateVec_7_state_valid <= _GEN_3027;
      end
    end else begin
      stateVec_7_state_valid <= _GEN_3027;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_7_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h7 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_7_state_inflight <= 1'h0;
      end else begin
        stateVec_7_state_inflight <= _GEN_3011;
      end
    end else begin
      stateVec_7_state_inflight <= _GEN_3011;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_7_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_7_w_timeout <= _GEN_3171; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h7 == sbuffer_out_s0_evictionIdx) begin
        stateVec_7_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_7_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_871) begin // @[Sbuffer.scala 745:8]
      stateVec_7_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_760) begin // @[Sbuffer.scala 511:20]
      stateVec_7_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_7_w_sameblock_inflight <= _GEN_314;
      end else begin
        stateVec_7_w_sameblock_inflight <= _GEN_457;
      end
    end else begin
      stateVec_7_w_sameblock_inflight <= _GEN_314;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_8_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h8 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_8_state_valid <= 1'h0;
      end else begin
        stateVec_8_state_valid <= _GEN_3028;
      end
    end else begin
      stateVec_8_state_valid <= _GEN_3028;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_8_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h8 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_8_state_inflight <= 1'h0;
      end else begin
        stateVec_8_state_inflight <= _GEN_3012;
      end
    end else begin
      stateVec_8_state_inflight <= _GEN_3012;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_8_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_8_w_timeout <= _GEN_3172; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h8 == sbuffer_out_s0_evictionIdx) begin
        stateVec_8_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_8_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_877) begin // @[Sbuffer.scala 745:8]
      stateVec_8_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_766) begin // @[Sbuffer.scala 511:20]
      stateVec_8_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_8_w_sameblock_inflight <= _GEN_319;
      end else begin
        stateVec_8_w_sameblock_inflight <= _GEN_464;
      end
    end else begin
      stateVec_8_w_sameblock_inflight <= _GEN_319;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_9_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h9 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_9_state_valid <= 1'h0;
      end else begin
        stateVec_9_state_valid <= _GEN_3029;
      end
    end else begin
      stateVec_9_state_valid <= _GEN_3029;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_9_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'h9 == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_9_state_inflight <= 1'h0;
      end else begin
        stateVec_9_state_inflight <= _GEN_3013;
      end
    end else begin
      stateVec_9_state_inflight <= _GEN_3013;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_9_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_9_w_timeout <= _GEN_3173; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'h9 == sbuffer_out_s0_evictionIdx) begin
        stateVec_9_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_9_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_883) begin // @[Sbuffer.scala 745:8]
      stateVec_9_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_772) begin // @[Sbuffer.scala 511:20]
      stateVec_9_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_9_w_sameblock_inflight <= _GEN_324;
      end else begin
        stateVec_9_w_sameblock_inflight <= _GEN_471;
      end
    end else begin
      stateVec_9_w_sameblock_inflight <= _GEN_324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_10_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'ha == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_10_state_valid <= 1'h0;
      end else begin
        stateVec_10_state_valid <= _GEN_3030;
      end
    end else begin
      stateVec_10_state_valid <= _GEN_3030;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_10_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'ha == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_10_state_inflight <= 1'h0;
      end else begin
        stateVec_10_state_inflight <= _GEN_3014;
      end
    end else begin
      stateVec_10_state_inflight <= _GEN_3014;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_10_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_10_w_timeout <= _GEN_3174; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'ha == sbuffer_out_s0_evictionIdx) begin
        stateVec_10_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_10_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_889) begin // @[Sbuffer.scala 745:8]
      stateVec_10_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_778) begin // @[Sbuffer.scala 511:20]
      stateVec_10_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_10_w_sameblock_inflight <= _GEN_329;
      end else begin
        stateVec_10_w_sameblock_inflight <= _GEN_478;
      end
    end else begin
      stateVec_10_w_sameblock_inflight <= _GEN_329;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_11_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hb == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_11_state_valid <= 1'h0;
      end else begin
        stateVec_11_state_valid <= _GEN_3031;
      end
    end else begin
      stateVec_11_state_valid <= _GEN_3031;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_11_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hb == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_11_state_inflight <= 1'h0;
      end else begin
        stateVec_11_state_inflight <= _GEN_3015;
      end
    end else begin
      stateVec_11_state_inflight <= _GEN_3015;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_11_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_11_w_timeout <= _GEN_3175; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'hb == sbuffer_out_s0_evictionIdx) begin
        stateVec_11_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_11_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_895) begin // @[Sbuffer.scala 745:8]
      stateVec_11_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_784) begin // @[Sbuffer.scala 511:20]
      stateVec_11_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_11_w_sameblock_inflight <= _GEN_334;
      end else begin
        stateVec_11_w_sameblock_inflight <= _GEN_485;
      end
    end else begin
      stateVec_11_w_sameblock_inflight <= _GEN_334;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_12_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hc == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_12_state_valid <= 1'h0;
      end else begin
        stateVec_12_state_valid <= _GEN_3032;
      end
    end else begin
      stateVec_12_state_valid <= _GEN_3032;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_12_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hc == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_12_state_inflight <= 1'h0;
      end else begin
        stateVec_12_state_inflight <= _GEN_3016;
      end
    end else begin
      stateVec_12_state_inflight <= _GEN_3016;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_12_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_12_w_timeout <= _GEN_3176; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'hc == sbuffer_out_s0_evictionIdx) begin
        stateVec_12_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_12_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_901) begin // @[Sbuffer.scala 745:8]
      stateVec_12_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_790) begin // @[Sbuffer.scala 511:20]
      stateVec_12_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_12_w_sameblock_inflight <= _GEN_339;
      end else begin
        stateVec_12_w_sameblock_inflight <= _GEN_492;
      end
    end else begin
      stateVec_12_w_sameblock_inflight <= _GEN_339;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_13_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hd == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_13_state_valid <= 1'h0;
      end else begin
        stateVec_13_state_valid <= _GEN_3033;
      end
    end else begin
      stateVec_13_state_valid <= _GEN_3033;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_13_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hd == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_13_state_inflight <= 1'h0;
      end else begin
        stateVec_13_state_inflight <= _GEN_3017;
      end
    end else begin
      stateVec_13_state_inflight <= _GEN_3017;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_13_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_13_w_timeout <= _GEN_3177; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'hd == sbuffer_out_s0_evictionIdx) begin
        stateVec_13_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_13_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_907) begin // @[Sbuffer.scala 745:8]
      stateVec_13_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_796) begin // @[Sbuffer.scala 511:20]
      stateVec_13_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_13_w_sameblock_inflight <= _GEN_344;
      end else begin
        stateVec_13_w_sameblock_inflight <= _GEN_499;
      end
    end else begin
      stateVec_13_w_sameblock_inflight <= _GEN_344;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_14_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'he == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_14_state_valid <= 1'h0;
      end else begin
        stateVec_14_state_valid <= _GEN_3034;
      end
    end else begin
      stateVec_14_state_valid <= _GEN_3034;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_14_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'he == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_14_state_inflight <= 1'h0;
      end else begin
        stateVec_14_state_inflight <= _GEN_3018;
      end
    end else begin
      stateVec_14_state_inflight <= _GEN_3018;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_14_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_14_w_timeout <= _GEN_3178; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'he == sbuffer_out_s0_evictionIdx) begin
        stateVec_14_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_14_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_913) begin // @[Sbuffer.scala 745:8]
      stateVec_14_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_802) begin // @[Sbuffer.scala 511:20]
      stateVec_14_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_14_w_sameblock_inflight <= _GEN_349;
      end else begin
        stateVec_14_w_sameblock_inflight <= _GEN_506;
      end
    end else begin
      stateVec_14_w_sameblock_inflight <= _GEN_349;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_15_state_valid <= 1'h0; // @[Sbuffer.scala 728:{44,44}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hf == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_15_state_valid <= 1'h0;
      end else begin
        stateVec_15_state_valid <= _GEN_3035;
      end
    end else begin
      stateVec_15_state_valid <= _GEN_3035;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 726:24]
      stateVec_15_state_inflight <= 1'h0; // @[Sbuffer.scala 727:{47,47}]
    end else if (io_dcache_refill_hit_resp_valid) begin
      if (4'hf == io_dcache_refill_hit_resp_bits_id[3:0]) begin
        stateVec_15_state_inflight <= 1'h0;
      end else begin
        stateVec_15_state_inflight <= _GEN_3019;
      end
    end else begin
      stateVec_15_state_inflight <= _GEN_3019;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 758:39]
      stateVec_15_w_timeout <= 1'h0;
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 678:28]
      stateVec_15_w_timeout <= _GEN_3179; // @[Sbuffer.scala 280:25 680:{52,52}]
    end else if (sbuffer_out_s0_fire) begin // @[Sbuffer.scala 280:25]
      if (4'hf == sbuffer_out_s0_evictionIdx) begin
        stateVec_15_w_timeout <= 1'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 745:8]
      stateVec_15_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_919) begin // @[Sbuffer.scala 745:8]
      stateVec_15_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 746:42]
    end else if (_T_808) begin // @[Sbuffer.scala 511:20]
      stateVec_15_w_sameblock_inflight <= 1'h0; // @[Sbuffer.scala 512:24]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        stateVec_15_w_sameblock_inflight <= _GEN_354;
      end else begin
        stateVec_15_w_sameblock_inflight <= _GEN_513;
      end
    end else begin
      stateVec_15_w_sameblock_inflight <= _GEN_354;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_0 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_1 & ~cohTimeOutMask_0) begin // @[Sbuffer.scala 511:20]
      cohCount_0 <= _cohCount_0_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[0]) begin
          cohCount_0 <= 21'h0;
        end else begin
          cohCount_0 <= _GEN_261;
        end
      end else if (secondInsertVec[0]) begin
        cohCount_0 <= 21'h0;
      end else begin
        cohCount_0 <= _GEN_261;
      end
    end else begin
      cohCount_0 <= _GEN_261;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_1 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_5 & ~cohTimeOutMask_1) begin // @[Sbuffer.scala 511:20]
      cohCount_1 <= _cohCount_1_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[1]) begin
          cohCount_1 <= 21'h0;
        end else begin
          cohCount_1 <= _GEN_263;
        end
      end else if (secondInsertVec[1]) begin
        cohCount_1 <= 21'h0;
      end else begin
        cohCount_1 <= _GEN_263;
      end
    end else begin
      cohCount_1 <= _GEN_263;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_2 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_9 & ~cohTimeOutMask_2) begin // @[Sbuffer.scala 511:20]
      cohCount_2 <= _cohCount_2_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[2]) begin
          cohCount_2 <= 21'h0;
        end else begin
          cohCount_2 <= _GEN_264;
        end
      end else if (secondInsertVec[2]) begin
        cohCount_2 <= 21'h0;
      end else begin
        cohCount_2 <= _GEN_264;
      end
    end else begin
      cohCount_2 <= _GEN_264;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_3 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_13 & ~cohTimeOutMask_3) begin // @[Sbuffer.scala 511:20]
      cohCount_3 <= _cohCount_3_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[3]) begin
          cohCount_3 <= 21'h0;
        end else begin
          cohCount_3 <= _GEN_265;
        end
      end else if (secondInsertVec[3]) begin
        cohCount_3 <= 21'h0;
      end else begin
        cohCount_3 <= _GEN_265;
      end
    end else begin
      cohCount_3 <= _GEN_265;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_4 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_17 & ~cohTimeOutMask_4) begin // @[Sbuffer.scala 511:20]
      cohCount_4 <= _cohCount_4_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[4]) begin
          cohCount_4 <= 21'h0;
        end else begin
          cohCount_4 <= _GEN_266;
        end
      end else if (secondInsertVec[4]) begin
        cohCount_4 <= 21'h0;
      end else begin
        cohCount_4 <= _GEN_266;
      end
    end else begin
      cohCount_4 <= _GEN_266;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_5 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_21 & ~cohTimeOutMask_5) begin // @[Sbuffer.scala 511:20]
      cohCount_5 <= _cohCount_5_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[5]) begin
          cohCount_5 <= 21'h0;
        end else begin
          cohCount_5 <= _GEN_267;
        end
      end else if (secondInsertVec[5]) begin
        cohCount_5 <= 21'h0;
      end else begin
        cohCount_5 <= _GEN_267;
      end
    end else begin
      cohCount_5 <= _GEN_267;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_6 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_25 & ~cohTimeOutMask_6) begin // @[Sbuffer.scala 511:20]
      cohCount_6 <= _cohCount_6_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[6]) begin
          cohCount_6 <= 21'h0;
        end else begin
          cohCount_6 <= _GEN_268;
        end
      end else if (secondInsertVec[6]) begin
        cohCount_6 <= 21'h0;
      end else begin
        cohCount_6 <= _GEN_268;
      end
    end else begin
      cohCount_6 <= _GEN_268;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_7 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_29 & ~cohTimeOutMask_7) begin // @[Sbuffer.scala 511:20]
      cohCount_7 <= _cohCount_7_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[7]) begin
          cohCount_7 <= 21'h0;
        end else begin
          cohCount_7 <= _GEN_269;
        end
      end else if (secondInsertVec[7]) begin
        cohCount_7 <= 21'h0;
      end else begin
        cohCount_7 <= _GEN_269;
      end
    end else begin
      cohCount_7 <= _GEN_269;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_8 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_33 & ~cohTimeOutMask_8) begin // @[Sbuffer.scala 511:20]
      cohCount_8 <= _cohCount_8_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[8]) begin
          cohCount_8 <= 21'h0;
        end else begin
          cohCount_8 <= _GEN_270;
        end
      end else if (secondInsertVec[8]) begin
        cohCount_8 <= 21'h0;
      end else begin
        cohCount_8 <= _GEN_270;
      end
    end else begin
      cohCount_8 <= _GEN_270;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_9 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_37 & ~cohTimeOutMask_9) begin // @[Sbuffer.scala 511:20]
      cohCount_9 <= _cohCount_9_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[9]) begin
          cohCount_9 <= 21'h0;
        end else begin
          cohCount_9 <= _GEN_271;
        end
      end else if (secondInsertVec[9]) begin
        cohCount_9 <= 21'h0;
      end else begin
        cohCount_9 <= _GEN_271;
      end
    end else begin
      cohCount_9 <= _GEN_271;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_10 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_41 & ~cohTimeOutMask_10) begin // @[Sbuffer.scala 511:20]
      cohCount_10 <= _cohCount_10_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[10]) begin
          cohCount_10 <= 21'h0;
        end else begin
          cohCount_10 <= _GEN_272;
        end
      end else if (secondInsertVec[10]) begin
        cohCount_10 <= 21'h0;
      end else begin
        cohCount_10 <= _GEN_272;
      end
    end else begin
      cohCount_10 <= _GEN_272;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_11 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_45 & ~cohTimeOutMask_11) begin // @[Sbuffer.scala 511:20]
      cohCount_11 <= _cohCount_11_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[11]) begin
          cohCount_11 <= 21'h0;
        end else begin
          cohCount_11 <= _GEN_273;
        end
      end else if (secondInsertVec[11]) begin
        cohCount_11 <= 21'h0;
      end else begin
        cohCount_11 <= _GEN_273;
      end
    end else begin
      cohCount_11 <= _GEN_273;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_12 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_49 & ~cohTimeOutMask_12) begin // @[Sbuffer.scala 511:20]
      cohCount_12 <= _cohCount_12_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[12]) begin
          cohCount_12 <= 21'h0;
        end else begin
          cohCount_12 <= _GEN_274;
        end
      end else if (secondInsertVec[12]) begin
        cohCount_12 <= 21'h0;
      end else begin
        cohCount_12 <= _GEN_274;
      end
    end else begin
      cohCount_12 <= _GEN_274;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_13 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_53 & ~cohTimeOutMask_13) begin // @[Sbuffer.scala 511:20]
      cohCount_13 <= _cohCount_13_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[13]) begin
          cohCount_13 <= 21'h0;
        end else begin
          cohCount_13 <= _GEN_275;
        end
      end else if (secondInsertVec[13]) begin
        cohCount_13 <= 21'h0;
      end else begin
        cohCount_13 <= _GEN_275;
      end
    end else begin
      cohCount_13 <= _GEN_275;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_14 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_57 & ~cohTimeOutMask_14) begin // @[Sbuffer.scala 511:20]
      cohCount_14 <= _cohCount_14_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[14]) begin
          cohCount_14 <= 21'h0;
        end else begin
          cohCount_14 <= _GEN_276;
        end
      end else if (secondInsertVec[14]) begin
        cohCount_14 <= 21'h0;
      end else begin
        cohCount_14 <= _GEN_276;
      end
    end else begin
      cohCount_14 <= _GEN_276;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 771:46]
      cohCount_15 <= 21'h0; // @[Sbuffer.scala 772:19]
    end else if (_candidateVec_T_61 & ~cohTimeOutMask_15) begin // @[Sbuffer.scala 511:20]
      cohCount_15 <= _cohCount_15_T_1; // @[Sbuffer.scala 512:24 482:32 483:28 458:32 464:28]
    end else if (_dataModule_io_writeReq_1_valid_T) begin
      if (canMerge_1) begin
        if (mergeVec_1[15]) begin
          cohCount_15 <= 21'h0;
        end else begin
          cohCount_15 <= _GEN_277;
        end
      end else if (secondInsertVec[15]) begin
        cohCount_15 <= 21'h0;
      end else begin
        cohCount_15 <= _GEN_277;
      end
    end else begin
      cohCount_15 <= _GEN_277;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_0 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_0_w_timeout & stateVec_0_state_inflight & ~missqReplayCount_0[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_0 <= _missqReplayCount_0_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h0 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_0 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_1 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_1_w_timeout & stateVec_1_state_inflight & ~missqReplayCount_1[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_1 <= _missqReplayCount_1_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h1 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_1 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_2 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_2_w_timeout & stateVec_2_state_inflight & ~missqReplayCount_2[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_2 <= _missqReplayCount_2_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h2 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_2 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_3 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_3_w_timeout & stateVec_3_state_inflight & ~missqReplayCount_3[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_3 <= _missqReplayCount_3_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h3 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_3 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_4 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_4_w_timeout & stateVec_4_state_inflight & ~missqReplayCount_4[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_4 <= _missqReplayCount_4_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h4 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_4 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_5 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_5_w_timeout & stateVec_5_state_inflight & ~missqReplayCount_5[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_5 <= _missqReplayCount_5_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h5 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_5 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_6 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_6_w_timeout & stateVec_6_state_inflight & ~missqReplayCount_6[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_6 <= _missqReplayCount_6_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h6 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_6 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_7 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_7_w_timeout & stateVec_7_state_inflight & ~missqReplayCount_7[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_7 <= _missqReplayCount_7_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h7 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_7 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_8 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_8_w_timeout & stateVec_8_state_inflight & ~missqReplayCount_8[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_8 <= _missqReplayCount_8_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h8 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_8 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_9 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_9_w_timeout & stateVec_9_state_inflight & ~missqReplayCount_9[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_9 <= _missqReplayCount_9_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'h9 == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_9 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_10 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_10_w_timeout & stateVec_10_state_inflight & ~missqReplayCount_10[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_10 <= _missqReplayCount_10_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'ha == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_10 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_11 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_11_w_timeout & stateVec_11_state_inflight & ~missqReplayCount_11[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_11 <= _missqReplayCount_11_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'hb == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_11 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_12 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_12_w_timeout & stateVec_12_state_inflight & ~missqReplayCount_12[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_12 <= _missqReplayCount_12_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'hc == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_12 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_13 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_13_w_timeout & stateVec_13_state_inflight & ~missqReplayCount_13[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_13 <= _missqReplayCount_13_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'hd == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_13 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_14 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_14_w_timeout & stateVec_14_state_inflight & ~missqReplayCount_14[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_14 <= _missqReplayCount_14_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'he == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_14 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 768:111]
      missqReplayCount_15 <= 5'h0; // @[Sbuffer.scala 769:27]
    end else if (stateVec_15_w_timeout & stateVec_15_state_inflight & ~missqReplayCount_15[4]) begin // @[Sbuffer.scala 758:39]
      missqReplayCount_15 <= _missqReplayCount_15_T_1; // @[Sbuffer.scala 282:33 759:{38,38}]
    end else if (io_dcache_replay_resp_valid) begin // @[Sbuffer.scala 282:33]
      if (4'hf == io_dcache_replay_resp_bits_id[3:0]) begin
        missqReplayCount_15 <= 5'h0;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 559:24]
      sbuffer_state <= 2'h0; // @[Sbuffer.scala 561:27 562:23 563:33 564:23 565:30 566:23 295:30]
    end else if (2'h0 == sbuffer_state) begin // @[Sbuffer.scala 559:24]
      if (io_flush_valid) begin // @[Sbuffer.scala 570:18]
        sbuffer_state <= 2'h2; // @[Sbuffer.scala 571:23]
      end else if (do_uarch_drain) begin // @[Sbuffer.scala 295:30]
        sbuffer_state <= 2'h3;
      end else if (do_eviction) begin
        sbuffer_state <= 2'h1;
      end
    end else if (2'h2 == sbuffer_state) begin // @[Sbuffer.scala 559:24]
      if (empty) begin // @[Sbuffer.scala 575:27]
        sbuffer_state <= 2'h0; // @[Sbuffer.scala 576:23]
      end
    end else if (2'h3 == sbuffer_state) begin // @[Sbuffer.scala 559:24]
      if (io_flush_valid) begin
        sbuffer_state <= 2'h2;
      end else begin
        sbuffer_state <= _GEN_718;
      end
    end else if (2'h1 == sbuffer_state) begin // @[Sbuffer.scala 295:30]
      sbuffer_state <= _GEN_722;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 420:24]
      enbufferSelReg <= 1'h0; // @[Sbuffer.scala 421:20]
    end else if (io_in_0_valid) begin // @[Sbuffer.scala 419:31]
      enbufferSelReg <= ~enbufferSelReg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 552:95]
      do_eviction <= 1'h0;
    end else begin
      do_eviction <= ActiveCount >= threshold | ActiveCount == 5'hf | ValidCount == 5'h10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 675:29]
      sbuffer_out_s1_valid <= 1'h0; // @[Sbuffer.scala 676:26]
    end else if (sbuffer_out_s0_cango) begin // @[Sbuffer.scala 671:28]
      sbuffer_out_s1_valid <= sbuffer_out_s0_valid; // @[Sbuffer.scala 672:26]
    end else if (sbuffer_out_s1_fire) begin // @[Sbuffer.scala 666:37]
      sbuffer_out_s1_valid <= 1'h0;
    end
  end
endmodule