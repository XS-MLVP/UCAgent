module bosc_Ifu(
  input          clock,
  input          reset,
  output         io_fromFtq_req_ready,
  input          io_fromFtq_req_valid,
  input          io_fromFtq_req_bits_fetch_0_valid,
  input  [48:0]  io_fromFtq_req_bits_fetch_0_startVAddr_addr,
  input  [48:0]  io_fromFtq_req_bits_fetch_0_nextStartVAddr_addr,
  input          io_fromFtq_req_bits_fetch_0_ftqIdx_flag,
  input  [5:0]   io_fromFtq_req_bits_fetch_0_ftqIdx_value,
  input          io_fromFtq_req_bits_fetch_0_takenCfiOffset_valid,
  input  [4:0]   io_fromFtq_req_bits_fetch_0_takenCfiOffset_bits,
  input          io_fromFtq_redirect_valid,
  input          io_fromFtq_flushFromBpu_s3_valid,
  input          io_fromFtq_flushFromBpu_s3_bits_flag,
  input  [5:0]   io_fromFtq_flushFromBpu_s3_bits_value,
  output         io_toFtq_wbRedirect_valid,
  output         io_toFtq_wbRedirect_bits_ftqIdx_flag,
  output [5:0]   io_toFtq_wbRedirect_bits_ftqIdx_value,
  output [49:0]  io_toFtq_wbRedirect_bits_pc,
  output         io_toFtq_wbRedirect_bits_taken,
  output [4:0]   io_toFtq_wbRedirect_bits_ftqOffset,
  output         io_toFtq_wbRedirect_bits_isRVC,
  output [1:0]   io_toFtq_wbRedirect_bits_attribute_rasAction,
  output [49:0]  io_toFtq_wbRedirect_bits_target,
  input          io_fromICache_fetchResp_valid,
  input          io_fromICache_fetchResp_bits_doubleline,
  input  [48:0]  io_fromICache_fetchResp_bits_vAddr_0_addr,
  input  [511:0] io_fromICache_fetchResp_bits_data,
  input  [31:0]  io_fromICache_fetchResp_bits_maybeRvcMap,
  input  [46:0]  io_fromICache_fetchResp_bits_pAddr_addr,
  input  [2:0]   io_fromICache_fetchResp_bits_exception_value,
  input          io_fromICache_fetchResp_bits_pmpMmio,
  input  [1:0]   io_fromICache_fetchResp_bits_itlbPbmt,
  input          io_fromICache_fetchResp_bits_isBackendException,
  input  [54:0]  io_fromICache_fetchResp_bits_gpAddr_addr,
  input          io_fromICache_fetchResp_bits_isForVSnonLeafPTE,
  input          io_fromICache_perf_hits_0,
  input          io_fromICache_perf_hits_1,
  input          io_fromICache_perf_isDoubleLine,
  input          io_fromICache_fetchReady,
  output         io_toICache_stall,
  input          io_toUncache_req_ready,
  output         io_toUncache_req_valid,
  output [46:0]  io_toUncache_req_bits_addr_addr,
  input          io_fromUncache_resp_valid,
  input  [31:0]  io_fromUncache_resp_bits_data,
  input          io_fromUncache_resp_bits_corrupt,
  input          io_fromUncache_resp_bits_denied,
  input          io_fromUncache_resp_bits_incomplete,
  input          io_toIBuffer_ready,
  output         io_toIBuffer_valid,
  output [31:0]  io_toIBuffer_bits_instrs_0,
  output [31:0]  io_toIBuffer_bits_instrs_1,
  output [31:0]  io_toIBuffer_bits_instrs_2,
  output [31:0]  io_toIBuffer_bits_instrs_3,
  output [31:0]  io_toIBuffer_bits_instrs_4,
  output [31:0]  io_toIBuffer_bits_instrs_5,
  output [31:0]  io_toIBuffer_bits_instrs_6,
  output [31:0]  io_toIBuffer_bits_instrs_7,
  output [31:0]  io_toIBuffer_bits_instrs_8,
  output [31:0]  io_toIBuffer_bits_instrs_9,
  output [31:0]  io_toIBuffer_bits_instrs_10,
  output [31:0]  io_toIBuffer_bits_instrs_11,
  output [31:0]  io_toIBuffer_bits_instrs_12,
  output [31:0]  io_toIBuffer_bits_instrs_13,
  output [31:0]  io_toIBuffer_bits_instrs_14,
  output [31:0]  io_toIBuffer_bits_instrs_15,
  output [31:0]  io_toIBuffer_bits_instrs_16,
  output [31:0]  io_toIBuffer_bits_instrs_17,
  output [31:0]  io_toIBuffer_bits_instrs_18,
  output [31:0]  io_toIBuffer_bits_instrs_19,
  output [31:0]  io_toIBuffer_bits_instrs_20,
  output [31:0]  io_toIBuffer_bits_instrs_21,
  output [31:0]  io_toIBuffer_bits_instrs_22,
  output [31:0]  io_toIBuffer_bits_instrs_23,
  output [31:0]  io_toIBuffer_bits_instrs_24,
  output [31:0]  io_toIBuffer_bits_instrs_25,
  output [31:0]  io_toIBuffer_bits_instrs_26,
  output [31:0]  io_toIBuffer_bits_instrs_27,
  output [31:0]  io_toIBuffer_bits_instrs_28,
  output [31:0]  io_toIBuffer_bits_instrs_29,
  output [31:0]  io_toIBuffer_bits_instrs_30,
  output [31:0]  io_toIBuffer_bits_instrs_31,
  output [31:0]  io_toIBuffer_bits_instrs_32,
  output [31:0]  io_toIBuffer_bits_instrs_33,
  output [31:0]  io_toIBuffer_bits_instrs_34,
  output [31:0]  io_toIBuffer_bits_instrs_35,
  output [35:0]  io_toIBuffer_bits_valid,
  output [35:0]  io_toIBuffer_bits_enqEnable,
  output         io_toIBuffer_bits_isRvc_0,
  output         io_toIBuffer_bits_isRvc_1,
  output         io_toIBuffer_bits_isRvc_2,
  output         io_toIBuffer_bits_isRvc_3,
  output         io_toIBuffer_bits_isRvc_4,
  output         io_toIBuffer_bits_isRvc_5,
  output         io_toIBuffer_bits_isRvc_6,
  output         io_toIBuffer_bits_isRvc_7,
  output         io_toIBuffer_bits_isRvc_8,
  output         io_toIBuffer_bits_isRvc_9,
  output         io_toIBuffer_bits_isRvc_10,
  output         io_toIBuffer_bits_isRvc_11,
  output         io_toIBuffer_bits_isRvc_12,
  output         io_toIBuffer_bits_isRvc_13,
  output         io_toIBuffer_bits_isRvc_14,
  output         io_toIBuffer_bits_isRvc_15,
  output         io_toIBuffer_bits_isRvc_16,
  output         io_toIBuffer_bits_isRvc_17,
  output         io_toIBuffer_bits_isRvc_18,
  output         io_toIBuffer_bits_isRvc_19,
  output         io_toIBuffer_bits_isRvc_20,
  output         io_toIBuffer_bits_isRvc_21,
  output         io_toIBuffer_bits_isRvc_22,
  output         io_toIBuffer_bits_isRvc_23,
  output         io_toIBuffer_bits_isRvc_24,
  output         io_toIBuffer_bits_isRvc_25,
  output         io_toIBuffer_bits_isRvc_26,
  output         io_toIBuffer_bits_isRvc_27,
  output         io_toIBuffer_bits_isRvc_28,
  output         io_toIBuffer_bits_isRvc_29,
  output         io_toIBuffer_bits_isRvc_30,
  output         io_toIBuffer_bits_isRvc_31,
  output         io_toIBuffer_bits_isRvc_32,
  output         io_toIBuffer_bits_isRvc_33,
  output         io_toIBuffer_bits_isRvc_34,
  output         io_toIBuffer_bits_isRvc_35,
  output         io_toIBuffer_bits_instrEndOffset_0_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_0_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_0_offset,
  output         io_toIBuffer_bits_instrEndOffset_1_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_1_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_1_offset,
  output         io_toIBuffer_bits_instrEndOffset_2_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_2_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_2_offset,
  output         io_toIBuffer_bits_instrEndOffset_3_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_3_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_3_offset,
  output         io_toIBuffer_bits_instrEndOffset_4_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_4_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_4_offset,
  output         io_toIBuffer_bits_instrEndOffset_5_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_5_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_5_offset,
  output         io_toIBuffer_bits_instrEndOffset_6_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_6_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_6_offset,
  output         io_toIBuffer_bits_instrEndOffset_7_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_7_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_7_offset,
  output         io_toIBuffer_bits_instrEndOffset_8_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_8_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_8_offset,
  output         io_toIBuffer_bits_instrEndOffset_9_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_9_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_9_offset,
  output         io_toIBuffer_bits_instrEndOffset_10_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_10_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_10_offset,
  output         io_toIBuffer_bits_instrEndOffset_11_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_11_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_11_offset,
  output         io_toIBuffer_bits_instrEndOffset_12_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_12_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_12_offset,
  output         io_toIBuffer_bits_instrEndOffset_13_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_13_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_13_offset,
  output         io_toIBuffer_bits_instrEndOffset_14_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_14_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_14_offset,
  output         io_toIBuffer_bits_instrEndOffset_15_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_15_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_15_offset,
  output         io_toIBuffer_bits_instrEndOffset_16_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_16_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_16_offset,
  output         io_toIBuffer_bits_instrEndOffset_17_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_17_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_17_offset,
  output         io_toIBuffer_bits_instrEndOffset_18_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_18_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_18_offset,
  output         io_toIBuffer_bits_instrEndOffset_19_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_19_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_19_offset,
  output         io_toIBuffer_bits_instrEndOffset_20_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_20_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_20_offset,
  output         io_toIBuffer_bits_instrEndOffset_21_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_21_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_21_offset,
  output         io_toIBuffer_bits_instrEndOffset_22_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_22_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_22_offset,
  output         io_toIBuffer_bits_instrEndOffset_23_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_23_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_23_offset,
  output         io_toIBuffer_bits_instrEndOffset_24_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_24_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_24_offset,
  output         io_toIBuffer_bits_instrEndOffset_25_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_25_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_25_offset,
  output         io_toIBuffer_bits_instrEndOffset_26_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_26_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_26_offset,
  output         io_toIBuffer_bits_instrEndOffset_27_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_27_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_27_offset,
  output         io_toIBuffer_bits_instrEndOffset_28_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_28_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_28_offset,
  output         io_toIBuffer_bits_instrEndOffset_29_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_29_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_29_offset,
  output         io_toIBuffer_bits_instrEndOffset_30_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_30_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_30_offset,
  output         io_toIBuffer_bits_instrEndOffset_31_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_31_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_31_offset,
  output         io_toIBuffer_bits_instrEndOffset_32_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_32_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_32_offset,
  output         io_toIBuffer_bits_instrEndOffset_33_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_33_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_33_offset,
  output         io_toIBuffer_bits_instrEndOffset_34_predTaken,
  output         io_toIBuffer_bits_instrEndOffset_34_fixedTaken,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_34_offset,
  output [4:0]   io_toIBuffer_bits_instrEndOffset_35_offset,
  output [2:0]   io_toIBuffer_bits_exceptionType_value,
  output         io_toIBuffer_bits_isBackendException,
  output         io_toIBuffer_bits_exceptionCrossPage,
  output [5:0]   io_toIBuffer_bits_exceptionOffset,
  output [3:0]   io_toIBuffer_bits_triggered_0,
  output [3:0]   io_toIBuffer_bits_triggered_1,
  output [3:0]   io_toIBuffer_bits_triggered_2,
  output [3:0]   io_toIBuffer_bits_triggered_3,
  output [3:0]   io_toIBuffer_bits_triggered_4,
  output [3:0]   io_toIBuffer_bits_triggered_5,
  output [3:0]   io_toIBuffer_bits_triggered_6,
  output [3:0]   io_toIBuffer_bits_triggered_7,
  output [3:0]   io_toIBuffer_bits_triggered_8,
  output [3:0]   io_toIBuffer_bits_triggered_9,
  output [3:0]   io_toIBuffer_bits_triggered_10,
  output [3:0]   io_toIBuffer_bits_triggered_11,
  output [3:0]   io_toIBuffer_bits_triggered_12,
  output [3:0]   io_toIBuffer_bits_triggered_13,
  output [3:0]   io_toIBuffer_bits_triggered_14,
  output [3:0]   io_toIBuffer_bits_triggered_15,
  output [3:0]   io_toIBuffer_bits_triggered_16,
  output [3:0]   io_toIBuffer_bits_triggered_17,
  output [3:0]   io_toIBuffer_bits_triggered_18,
  output [3:0]   io_toIBuffer_bits_triggered_19,
  output [3:0]   io_toIBuffer_bits_triggered_20,
  output [3:0]   io_toIBuffer_bits_triggered_21,
  output [3:0]   io_toIBuffer_bits_triggered_22,
  output [3:0]   io_toIBuffer_bits_triggered_23,
  output [3:0]   io_toIBuffer_bits_triggered_24,
  output [3:0]   io_toIBuffer_bits_triggered_25,
  output [3:0]   io_toIBuffer_bits_triggered_26,
  output [3:0]   io_toIBuffer_bits_triggered_27,
  output [3:0]   io_toIBuffer_bits_triggered_28,
  output [3:0]   io_toIBuffer_bits_triggered_29,
  output [3:0]   io_toIBuffer_bits_triggered_30,
  output [3:0]   io_toIBuffer_bits_triggered_31,
  output [3:0]   io_toIBuffer_bits_triggered_32,
  output [3:0]   io_toIBuffer_bits_triggered_33,
  output [3:0]   io_toIBuffer_bits_triggered_34,
  output [3:0]   io_toIBuffer_bits_triggered_35,
  output         io_toIBuffer_bits_isLastInFtqEntry_0,
  output         io_toIBuffer_bits_isLastInFtqEntry_1,
  output         io_toIBuffer_bits_isLastInFtqEntry_2,
  output         io_toIBuffer_bits_isLastInFtqEntry_3,
  output         io_toIBuffer_bits_isLastInFtqEntry_4,
  output         io_toIBuffer_bits_isLastInFtqEntry_5,
  output         io_toIBuffer_bits_isLastInFtqEntry_6,
  output         io_toIBuffer_bits_isLastInFtqEntry_7,
  output         io_toIBuffer_bits_isLastInFtqEntry_8,
  output         io_toIBuffer_bits_isLastInFtqEntry_9,
  output         io_toIBuffer_bits_isLastInFtqEntry_10,
  output         io_toIBuffer_bits_isLastInFtqEntry_11,
  output         io_toIBuffer_bits_isLastInFtqEntry_12,
  output         io_toIBuffer_bits_isLastInFtqEntry_13,
  output         io_toIBuffer_bits_isLastInFtqEntry_14,
  output         io_toIBuffer_bits_isLastInFtqEntry_15,
  output         io_toIBuffer_bits_isLastInFtqEntry_16,
  output         io_toIBuffer_bits_isLastInFtqEntry_17,
  output         io_toIBuffer_bits_isLastInFtqEntry_18,
  output         io_toIBuffer_bits_isLastInFtqEntry_19,
  output         io_toIBuffer_bits_isLastInFtqEntry_20,
  output         io_toIBuffer_bits_isLastInFtqEntry_21,
  output         io_toIBuffer_bits_isLastInFtqEntry_22,
  output         io_toIBuffer_bits_isLastInFtqEntry_23,
  output         io_toIBuffer_bits_isLastInFtqEntry_24,
  output         io_toIBuffer_bits_isLastInFtqEntry_25,
  output         io_toIBuffer_bits_isLastInFtqEntry_26,
  output         io_toIBuffer_bits_isLastInFtqEntry_27,
  output         io_toIBuffer_bits_isLastInFtqEntry_28,
  output         io_toIBuffer_bits_isLastInFtqEntry_29,
  output         io_toIBuffer_bits_isLastInFtqEntry_30,
  output         io_toIBuffer_bits_isLastInFtqEntry_31,
  output         io_toIBuffer_bits_isLastInFtqEntry_32,
  output         io_toIBuffer_bits_isLastInFtqEntry_33,
  output         io_toIBuffer_bits_isLastInFtqEntry_34,
  output         io_toIBuffer_bits_isLastInFtqEntry_35,
  output [48:0]  io_toIBuffer_bits_pc_0_addr,
  output [48:0]  io_toIBuffer_bits_pc_1_addr,
  output [48:0]  io_toIBuffer_bits_pc_2_addr,
  output [48:0]  io_toIBuffer_bits_pc_3_addr,
  output [48:0]  io_toIBuffer_bits_pc_4_addr,
  output [48:0]  io_toIBuffer_bits_pc_5_addr,
  output [48:0]  io_toIBuffer_bits_pc_6_addr,
  output [48:0]  io_toIBuffer_bits_pc_7_addr,
  output [48:0]  io_toIBuffer_bits_pc_8_addr,
  output [48:0]  io_toIBuffer_bits_pc_9_addr,
  output [48:0]  io_toIBuffer_bits_pc_10_addr,
  output [48:0]  io_toIBuffer_bits_pc_11_addr,
  output [48:0]  io_toIBuffer_bits_pc_12_addr,
  output [48:0]  io_toIBuffer_bits_pc_13_addr,
  output [48:0]  io_toIBuffer_bits_pc_14_addr,
  output [48:0]  io_toIBuffer_bits_pc_15_addr,
  output [48:0]  io_toIBuffer_bits_pc_16_addr,
  output [48:0]  io_toIBuffer_bits_pc_17_addr,
  output [48:0]  io_toIBuffer_bits_pc_18_addr,
  output [48:0]  io_toIBuffer_bits_pc_19_addr,
  output [48:0]  io_toIBuffer_bits_pc_20_addr,
  output [48:0]  io_toIBuffer_bits_pc_21_addr,
  output [48:0]  io_toIBuffer_bits_pc_22_addr,
  output [48:0]  io_toIBuffer_bits_pc_23_addr,
  output [48:0]  io_toIBuffer_bits_pc_24_addr,
  output [48:0]  io_toIBuffer_bits_pc_25_addr,
  output [48:0]  io_toIBuffer_bits_pc_26_addr,
  output [48:0]  io_toIBuffer_bits_pc_27_addr,
  output [48:0]  io_toIBuffer_bits_pc_28_addr,
  output [48:0]  io_toIBuffer_bits_pc_29_addr,
  output [48:0]  io_toIBuffer_bits_pc_30_addr,
  output [48:0]  io_toIBuffer_bits_pc_31_addr,
  output [48:0]  io_toIBuffer_bits_pc_32_addr,
  output [48:0]  io_toIBuffer_bits_pc_33_addr,
  output [48:0]  io_toIBuffer_bits_pc_34_addr,
  output [48:0]  io_toIBuffer_bits_pc_35_addr,
  output [5:0]   io_toIBuffer_bits_prevInstrCount,
  output         io_toIBuffer_bits_ftqPtr_0_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_0_value,
  output         io_toIBuffer_bits_ftqPtr_1_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_1_value,
  output         io_toIBuffer_bits_ftqPtr_2_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_2_value,
  output         io_toIBuffer_bits_ftqPtr_3_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_3_value,
  output         io_toIBuffer_bits_ftqPtr_4_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_4_value,
  output         io_toIBuffer_bits_ftqPtr_5_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_5_value,
  output         io_toIBuffer_bits_ftqPtr_6_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_6_value,
  output         io_toIBuffer_bits_ftqPtr_7_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_7_value,
  output         io_toIBuffer_bits_ftqPtr_8_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_8_value,
  output         io_toIBuffer_bits_ftqPtr_9_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_9_value,
  output         io_toIBuffer_bits_ftqPtr_10_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_10_value,
  output         io_toIBuffer_bits_ftqPtr_11_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_11_value,
  output         io_toIBuffer_bits_ftqPtr_12_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_12_value,
  output         io_toIBuffer_bits_ftqPtr_13_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_13_value,
  output         io_toIBuffer_bits_ftqPtr_14_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_14_value,
  output         io_toIBuffer_bits_ftqPtr_15_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_15_value,
  output         io_toIBuffer_bits_ftqPtr_16_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_16_value,
  output         io_toIBuffer_bits_ftqPtr_17_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_17_value,
  output         io_toIBuffer_bits_ftqPtr_18_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_18_value,
  output         io_toIBuffer_bits_ftqPtr_19_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_19_value,
  output         io_toIBuffer_bits_ftqPtr_20_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_20_value,
  output         io_toIBuffer_bits_ftqPtr_21_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_21_value,
  output         io_toIBuffer_bits_ftqPtr_22_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_22_value,
  output         io_toIBuffer_bits_ftqPtr_23_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_23_value,
  output         io_toIBuffer_bits_ftqPtr_24_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_24_value,
  output         io_toIBuffer_bits_ftqPtr_25_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_25_value,
  output         io_toIBuffer_bits_ftqPtr_26_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_26_value,
  output         io_toIBuffer_bits_ftqPtr_27_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_27_value,
  output         io_toIBuffer_bits_ftqPtr_28_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_28_value,
  output         io_toIBuffer_bits_ftqPtr_29_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_29_value,
  output         io_toIBuffer_bits_ftqPtr_30_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_30_value,
  output         io_toIBuffer_bits_ftqPtr_31_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_31_value,
  output         io_toIBuffer_bits_ftqPtr_32_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_32_value,
  output         io_toIBuffer_bits_ftqPtr_33_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_33_value,
  output         io_toIBuffer_bits_ftqPtr_34_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_34_value,
  output         io_toIBuffer_bits_ftqPtr_35_flag,
  output [5:0]   io_toIBuffer_bits_ftqPtr_35_value,
  output         io_toBackend_gpAddrMem_wen,
  output [5:0]   io_toBackend_gpAddrMem_waddr,
  output [55:0]  io_toBackend_gpAddrMem_wdata_gpaddr,
  output         io_toBackend_gpAddrMem_wdata_isForVSnonLeafPTE,
  input          io_frontendTrigger_tUpdate_valid,
  input  [1:0]   io_frontendTrigger_tUpdate_bits_addr,
  input  [1:0]   io_frontendTrigger_tUpdate_bits_tdata_matchType,
  input          io_frontendTrigger_tUpdate_bits_tdata_select,
  input  [3:0]   io_frontendTrigger_tUpdate_bits_tdata_action,
  input          io_frontendTrigger_tUpdate_bits_tdata_chain,
  input  [63:0]  io_frontendTrigger_tUpdate_bits_tdata_tdata2,
  input          io_frontendTrigger_tEnableVec_0,
  input          io_frontendTrigger_tEnableVec_1,
  input          io_frontendTrigger_tEnableVec_2,
  input          io_frontendTrigger_tEnableVec_3,
  input          io_frontendTrigger_debugMode,
  input          io_frontendTrigger_triggerCanRaiseBpExp,
  input          io_csrFsIsOff,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value,
  output [5:0]   io_perf_8_value,
  output [5:0]   io_perf_9_value,
  output [5:0]   io_perf_10_value,
  output [5:0]   io_perf_11_value,
  output [5:0]   io_perf_12_value
);

endmodule

